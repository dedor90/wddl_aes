
module aes_sbox_wddl ( a, a_n, d, d_n );
 input [7:0] a;
 input [7:0] a_n;
 output [7:0] d;
 output [7:0] d_n;
 wire  n2519, n2519_n, n2520, n2520_n, n2521, n2521_n, n2522, n2522_n, n2523, n2523_n, n2524, n2524_n, n2525, n2525_n, n2526, n2526_n, n2527, n2527_n, n2528, n2528_n, 
 n2529_n, n2529, n2530_n, n2530, n2531_n, n2531, n2532_n, n2532, n2533_n, n2533, n2534_n, n2534, n2535_n, n2535, n2536_n, n2536, n2537_n, n2537, n2538_n, n2538,
 n2539_n, n2539, n2540_n, n2540, n2541_n, n2541, n2542_n, n2542, n2543_n, n2543, n2544_n, n2544, n2545_n, n2545, n2546_n, n2546, n2547_n, n2547, n2548_n, n2548,
 n2549_n, n2549, n2550_n, n2550, n2551_n, n2551, n2552_n, n2552, n2553_n, n2553, n2554_n, n2554, n2555_n, n2555, n2556_n, n2556, n2557_n, n2557, n2558_n, n2558,
 n2559_n, n2559, n2560_n, n2560, n2561_n, n2561, n2562_n, n2562, n2563_n, n2563, n2564_n, n2564, n2565_n, n2565, n2566_n, n2566, n2567_n, n2567, n2568_n, n2568,
 n2569_n, n2569, n2570_n, n2570, n2571_n, n2571, n2572_n, n2572, n2573_n, n2573, n2574_n, n2574, n2575_n, n2575, n2576_n, n2576, n2577_n, n2577, n2578_n, n2578,
 n2579_n, n2579, n2580_n, n2580, n2581_n, n2581, n2582_n, n2582, n2583_n, n2583, n2584_n, n2584, n2585_n, n2585, n2586_n, n2586, n2587_n, n2587, n2588_n, n2588,
 n2589_n, n2589, n2590_n, n2590, n2591_n, n2591, n2592_n, n2592, n2593_n, n2593, n2594_n, n2594, n2595_n, n2595, n2596_n, n2596, n2597_n, n2597, n2598_n, n2598,
 n2599_n, n2599, n2600_n, n2600, n2601_n, n2601, n2602_n, n2602, n2603_n, n2603, n2604_n, n2604, n2605_n, n2605, n2606_n, n2606, n2607_n, n2607, n2608_n, n2608,
 n2609_n, n2609, n2610_n, n2610, n2611_n, n2611, n2612_n, n2612, n2613_n, n2613, n2614_n, n2614, n2615_n, n2615, n2616_n, n2616, n2617_n, n2617, n2618_n, n2618,
 n2619_n, n2619, n2620_n, n2620, n2621_n, n2621, n2622_n, n2622, n2623_n, n2623, n2624_n, n2624, n2625_n, n2625, n2626_n, n2626, n2627_n, n2627, n2628_n, n2628,
 n2629_n, n2629, n2630_n, n2630, n2631_n, n2631, n2632_n, n2632, n2633_n, n2633, n2634_n, n2634, n2635_n, n2635, n2636_n, n2636, n2637_n, n2637, n2638_n, n2638,
 n2639_n, n2639, n2640_n, n2640, n2641_n, n2641, n2642_n, n2642, n2643_n, n2643, n2644_n, n2644, n2645_n, n2645, n2646_n, n2646, n2647_n, n2647, n2648_n, n2648,
 n2649_n, n2649, n2650_n, n2650, n2651_n, n2651, n2652_n, n2652, n2653_n, n2653, n2654_n, n2654, n2655_n, n2655, n2656_n, n2656, n2657_n, n2657, n2658_n, n2658,
 n2659_n, n2659, n2660_n, n2660, n2661_n, n2661, n2662_n, n2662, n2663_n, n2663, n2664_n, n2664, n2665_n, n2665, n2666_n, n2666, n2667_n, n2667, n2668_n, n2668,
 n2669_n, n2669, n2670_n, n2670, n2671_n, n2671, n2672_n, n2672, n2673_n, n2673, n2674_n, n2674, n2675_n, n2675, n2676_n, n2676, n2677_n, n2677, n2678_n, n2678,
 n2679_n, n2679, n2680_n, n2680, n2681_n, n2681, n2682_n, n2682, n2683_n, n2683, n2684_n, n2684, n2685_n, n2685, n2686_n, n2686, n2687_n, n2687, n2688_n, n2688,
 n2689_n, n2689, n2690_n, n2690, n2691_n, n2691, n2692_n, n2692, n2693_n, n2693, n2694_n, n2694, n2695_n, n2695, n2696_n, n2696, n2697_n, n2697, n2698_n, n2698,
 n2699_n, n2699, n2700_n, n2700, n2701_n, n2701, n2702_n, n2702, n2703_n, n2703, n2704_n, n2704, n2705_n, n2705, n2706_n, n2706, n2707_n, n2707, n2708_n, n2708,
 n2709_n, n2709, n2710_n, n2710, n2711_n, n2711, n2712_n, n2712, n2713_n, n2713, n2714_n, n2714, n2715_n, n2715, n2716_n, n2716, n2717_n, n2717, n2718_n, n2718,
 n2719_n, n2719, n2720_n, n2720, n2721_n, n2721, n2722_n, n2722, n2723_n, n2723, n2724_n, n2724, n2725_n, n2725, n2726_n, n2726, n2727_n, n2727, n2728_n, n2728,
 n2729_n, n2729, n2730_n, n2730, n2731_n, n2731, n2732_n, n2732, n2733_n, n2733, n2734_n, n2734, n2735_n, n2735, n2736_n, n2736, n2737_n, n2737, n2738_n, n2738,
 n2739_n, n2739, n2740_n, n2740, n2741_n, n2741, n2742_n, n2742, n2743_n, n2743, n2744_n, n2744, n2745_n, n2745, n2746_n, n2746, n2747_n, n2747, n2748_n, n2748,
 n2749_n, n2749, n2750_n, n2750, n2751_n, n2751, n2752_n, n2752, n2753_n, n2753, n2754_n, n2754, n2755_n, n2755, n2756_n, n2756, n2757_n, n2757, n2758_n, n2758,
 n2759_n, n2759, n2760_n, n2760, n2761_n, n2761, n2762_n, n2762, n2763_n, n2763, n2764_n, n2764, n2765_n, n2765, n2766_n, n2766, n2767_n, n2767, n2768_n, n2768,
 n2769_n, n2769, n2770_n, n2770, n2771_n, n2771, n2772_n, n2772, n2773_n, n2773, n2774_n, n2774, n2775_n, n2775, n2776_n, n2776, n2777_n, n2777, n2778_n, n2778,
 n2779_n, n2779, n2780_n, n2780, n2781_n, n2781, n2782_n, n2782, n2783_n, n2783, n2784_n, n2784, n2785_n, n2785, n2786_n, n2786, n2787_n, n2787, n2788_n, n2788,
 n2789_n, n2789, n2790_n, n2790, n2791_n, n2791, n2792_n, n2792, n2793_n, n2793, n2794_n, n2794, n2795_n, n2795, n2796_n, n2796, n2797_n, n2797, n2798_n, n2798,
 n2799_n, n2799, n2800_n, n2800, n2801_n, n2801, n2802_n, n2802, n2803_n, n2803, n2804_n, n2804, n2805_n, n2805, n2806_n, n2806, n2807_n, n2807, n2808_n, n2808,
 n2809_n, n2809, n2810_n, n2810, n2811_n, n2811, n2812_n, n2812, n2813_n, n2813, n2814_n, n2814, n2815_n, n2815, n2816_n, n2816, n2817_n, n2817, n2818_n, n2818,
 n2819_n, n2819, n2820_n, n2820, n2821_n, n2821, n2822_n, n2822, n2823_n, n2823, n2824_n, n2824, n2825_n, n2825, n2826_n, n2826, n2827_n, n2827, n2828_n, n2828,
 n2829_n, n2829, n2830_n, n2830, n2831_n, n2831, n2832_n, n2832, n2833_n, n2833, n2834_n, n2834, n2835_n, n2835, n2836_n, n2836, n2837_n, n2837, n2838_n, n2838,
 n2839_n, n2839, n2840_n, n2840, n2841_n, n2841, n2842_n, n2842, n2843_n, n2843, n2844_n, n2844, n2845_n, n2845, n2846_n, n2846, n2847_n, n2847, n2848_n, n2848,
 n2849_n, n2849, n2850_n, n2850, n2851_n, n2851, n2852_n, n2852, n2853_n, n2853, n2854_n, n2854, n2855_n, n2855, n2856_n, n2856, n2857_n, n2857, n2858_n, n2858,
 n2859_n, n2859, n2860_n, n2860, n2861_n, n2861, n2862_n, n2862, n2863_n, n2863, n2864_n, n2864, n2865_n, n2865, n2866_n, n2866, n2867_n, n2867, n2868_n, n2868,
 n2869_n, n2869, n2870_n, n2870, n2871_n, n2871, n2872_n, n2872, n2873_n, n2873, n2874_n, n2874, n2875_n, n2875, n2876_n, n2876, n2877_n, n2877, n2878_n, n2878,
 n2879_n, n2879, n2880_n, n2880, n2881_n, n2881, n2882_n, n2882, n2883_n, n2883, n2884_n, n2884, n2885_n, n2885, n2886_n, n2886, n2887_n, n2887, n2888_n, n2888,
 n2889_n, n2889, n2890_n, n2890, n2891_n, n2891, n2892_n, n2892, n2893_n, n2893, n2894_n, n2894, n2895_n, n2895, n2896_n, n2896, n2897_n, n2897, n2898_n, n2898,
 n2899_n, n2899, n2900_n, n2900, n2901_n, n2901, n2902_n, n2902, n2903_n, n2903, n2904_n, n2904, n2905_n, n2905, n2906_n, n2906, n2907_n, n2907, n2908_n, n2908,
 n2909_n, n2909, n2910_n, n2910, n2911_n, n2911, n2912_n, n2912, n2913_n, n2913, n2914_n, n2914, n2915_n, n2915, n2916_n, n2916, n2917_n, n2917, n2918_n, n2918,
 n2919_n, n2919, n2920_n, n2920, n2921_n, n2921, n2922_n, n2922, n2923_n, n2923, n2924_n, n2924, n2925_n, n2925, n2926_n, n2926, n2927_n, n2927, n2928_n, n2928,
 n2929_n, n2929, n2930_n, n2930, n2931_n, n2931, n2932_n, n2932, n2933_n, n2933, n2934_n, n2934, n2935_n, n2935, n2936_n, n2936, n2937_n, n2937, n2938_n, n2938,
 n2939_n, n2939, n2940_n, n2940, n2941_n, n2941, n2942_n, n2942, n2943_n, n2943, n2944_n, n2944, n2945_n, n2945, n2946_n, n2946, n2947_n, n2947, n2948_n, n2948,
 n2949_n, n2949, n2950_n, n2950, n2951_n, n2951, n2952_n, n2952, n2953_n, n2953, n2954_n, n2954, n2955_n, n2955, n2956_n, n2956, n2957_n, n2957, n2958_n, n2958,
 n2959_n, n2959, n2960_n, n2960, n2961_n, n2961, n2962_n, n2962, n2963_n, n2963, n2964_n, n2964, n2965_n, n2965, n2966_n, n2966, n2967_n, n2967, n2968_n, n2968,
 n2969_n, n2969, n2970_n, n2970, n2971_n, n2971, n2972_n, n2972, n2973_n, n2973, n2974_n, n2974, n2975_n, n2975, n2976_n, n2976, n2977_n, n2977, n2978_n, n2978,
 n2979_n, n2979, n2980_n, n2980, n2981_n, n2981, n2982_n, n2982, n2983_n, n2983, n2984_n, n2984, n2985_n, n2985, n2986_n, n2986, n2987_n, n2987, n2988_n, n2988,
 n2989_n, n2989, n2990_n, n2990, n2991_n, n2991, n2992_n, n2992, n2993_n, n2993, n2994_n, n2994, n2995_n, n2995, n2996_n, n2996, n2997_n, n2997, n2998_n, n2998,
 n2999_n, n2999, n3000_n, n3000, n3001_n, n3001, n3002_n, n3002, n3003_n, n3003, n3004_n, n3004, n3005_n, n3005, n3006_n, n3006, n3007_n, n3007, n3008_n, n3008,
 n3009_n, n3009, n3010_n, n3010, n3011_n, n3011, n3012_n, n3012, n3013_n, n3013, n3014_n, n3014, n3015_n, n3015, n3016_n, n3016, n3017_n, n3017, n3018_n, n3018,
 n3019_n, n3019, n3020_n, n3020, n3021_n, n3021, n3022_n, n3022, n3023_n, n3023, n3024_n, n3024, n3025_n, n3025, n3026_n, n3026, n3027_n, n3027, n3028_n, n3028,
 n3029_n, n3029, n3030_n, n3030, n3031_n, n3031, n3032_n, n3032, n3033_n, n3033, n3034_n, n3034, n3035_n, n3035, n3036_n, n3036, n3037_n, n3037, n3038_n, n3038,
 n3039_n, n3039, n3040_n, n3040, n3041_n, n3041, n3042_n, n3042, n3043_n, n3043, n3044_n, n3044, n3045_n, n3045, n3046_n, n3046, n3047_n, n3047, n3048_n, n3048,
 n3049_n, n3049, n3050_n, n3050, n3051_n, n3051, n3052_n, n3052, n3053_n, n3053, n3054_n, n3054, n3055_n, n3055, n3056_n, n3056, n3057_n, n3057, n3058_n, n3058,
 n3059_n, n3059, n3060_n, n3060, n3061_n, n3061, n3062_n, n3062, n3063_n, n3063, n3064_n, n3064, n3065_n, n3065, n3066_n, n3066, n3067_n, n3067, n3068_n, n3068,
 n3069_n, n3069, n3070_n, n3070, n3071_n, n3071, n3072_n, n3072, n3073_n, n3073, n3074_n, n3074, n3075_n, n3075, n3076_n, n3076, n3077_n, n3077, n3078_n, n3078,
 n3079_n, n3079, n3080_n, n3080, n3081_n, n3081, n3082_n, n3082, n3083_n, n3083, n3084_n, n3084, n3085_n, n3085, n3086_n, n3086, n3087_n, n3087, n3088_n, n3088,
 n3089_n, n3089, n3090_n, n3090, n3091_n, n3091, n3092_n, n3092, n3093_n, n3093, n3094_n, n3094, n3095_n, n3095, n3096_n, n3096, n3097_n, n3097, n3098_n, n3098,
 n3099_n, n3099, n3100_n, n3100, n3101_n, n3101, n3102_n, n3102, n3103_n, n3103, n3104_n, n3104, n3105_n, n3105, n3106_n, n3106, n3107_n, n3107, n3108_n, n3108,
 n3109_n, n3109, n3110_n, n3110, n3111_n, n3111, n3112_n, n3112, n3113_n, n3113, n3114_n, n3114, n3115_n, n3115, n3116_n, n3116, n3117_n, n3117, n3118_n, n3118,
 n3119_n, n3119, n3120_n, n3120, n3121_n, n3121, n3122_n, n3122, n3123_n, n3123, n3124_n, n3124, n3125_n, n3125, n3126_n, n3126, n3127_n, n3127, n3128_n, n3128,
 n3129_n, n3129, n3130_n, n3130, n3131_n, n3131, n3132_n, n3132, n3133_n, n3133, n3134_n, n3134, n3135_n, n3135, n3136_n, n3136, n3137_n, n3137, n3138_n, n3138,
 n3139_n, n3139, n3140_n, n3140, n3141_n, n3141, n3142_n, n3142, n3143_n, n3143, n3144_n, n3144, n3145_n, n3145, n3146_n, n3146, n3147_n, n3147, n3148_n, n3148,
 n3149_n, n3149, n3150_n, n3150, n3151_n, n3151, n3152_n, n3152, n3153_n, n3153, n3154_n, n3154, n3155_n, n3155, n3156_n, n3156, n3157_n, n3157, n3158_n, n3158,
 n3159_n, n3159, n3160_n, n3160, n3161_n, n3161, n3162_n, n3162, n3163_n, n3163, n3164_n, n3164, n3165_n, n3165, n3166_n, n3166, n3167_n, n3167, n3168_n, n3168,
 n3169_n, n3169, n3170_n, n3170, n3171_n, n3171, n3172_n, n3172, n3173_n, n3173, n3174_n, n3174, n3175_n, n3175, n3176_n, n3176, n3177_n, n3177, n3178_n, n3178,
 n3179_n, n3179, n3180_n, n3180, n3181_n, n3181, n3182_n, n3182, n3183_n, n3183, n3184_n, n3184, n3185_n, n3185, n3186_n, n3186, n3187_n, n3187, n3188_n, n3188,
 n3189_n, n3189, n3190_n, n3190, n3191_n, n3191, n3192_n, n3192, n3193_n, n3193, n3194_n, n3194, n3195_n, n3195, n3196_n, n3196, n3197_n, n3197, n3198_n, n3198,
 n3199_n, n3199, n3200_n, n3200, n3201_n, n3201, n3202_n, n3202, n3203_n, n3203, n3204_n, n3204, n3205_n, n3205, n3206_n, n3206, n3207_n, n3207, n3208_n, n3208,
 n3209_n, n3209, n3210_n, n3210, n3211_n, n3211, n3212_n, n3212, n3213_n, n3213, n3214_n, n3214, n3215_n, n3215, n3216_n, n3216, n3217_n, n3217, n3218_n, n3218,
 n3219_n, n3219, n3220_n, n3220, n3221_n, n3221, n3222_n, n3222, n3223_n, n3223, n3224_n, n3224, n3225_n, n3225, n3226_n, n3226, n3227_n, n3227, n3228_n, n3228,
 n3229_n, n3229, n3230_n, n3230, n3231_n, n3231, n3232_n, n3232, n3233_n, n3233, n3234_n, n3234, n3235_n, n3235, n3236_n, n3236, n3237_n, n3237, n3238_n, n3238,
 n3239_n, n3239, n3240_n, n3240, n3241_n, n3241, n3242_n, n3242, n3243_n, n3243, n3244_n, n3244, n3245_n, n3245, n3246_n, n3246, n3247_n, n3247, n3248_n, n3248,
 n3249_n, n3249, n3250_n, n3250, n3251_n, n3251, n3252_n, n3252, n3253_n, n3253, n3254_n, n3254, n3255_n, n3255, n3256_n, n3256, n3257_n, n3257, n3258_n, n3258,
 n3259_n, n3259, n3260_n, n3260, n3261_n, n3261, n3262_n, n3262, n3263_n, n3263, n3264_n, n3264, n3265_n, n3265, n3266_n, n3266, n3267_n, n3267, n3268_n, n3268,
 n3269_n, n3269, n3270_n, n3270, n3271_n, n3271, n3272_n, n3272, n3273_n, n3273, n3274_n, n3274, n3275_n, n3275, n3276_n, n3276, n3277_n, n3277, n3278_n, n3278,
 n3279_n, n3279, n3280_n, n3280, n3281_n, n3281, n3282_n, n3282, n3283_n, n3283, n3284_n, n3284, n3285_n, n3285, n3286_n, n3286, n3287_n, n3287, n3288_n, n3288,
 n3289_n, n3289, n3290_n, n3290, n3291_n, n3291, n3292_n, n3292, n3293_n, n3293, n3294_n, n3294, n3295_n, n3295, n3296_n, n3296, n3297_n, n3297, n3298_n, n3298,
 n3299_n, n3299, n3300_n, n3300, n3301_n, n3301, n3302_n, n3302, n3303_n, n3303, n3304_n, n3304, n3305_n, n3305, n3306_n, n3306, n3307_n, n3307, n3308_n, n3308,
 n3309_n, n3309, n3310_n, n3310, n3311_n, n3311, n3312_n, n3312, n3313_n, n3313, n3314_n, n3314, n3315_n, n3315, n3316_n, n3316, n3317_n, n3317, n3318_n, n3318,
 n3319_n, n3319, n3320_n, n3320, n3321_n, n3321, n3322_n, n3322, n3323_n, n3323, n3324_n, n3324, n3325_n, n3325, n3326_n, n3326, n3327_n, n3327, n3328_n, n3328,
 n3329_n, n3329, n3330_n, n3330, n3331_n, n3331, n3332_n, n3332, n3333_n, n3333, n3334_n, n3334, n3335_n, n3335, n3336_n, n3336, n3337_n, n3337, n3338_n, n3338,
 n3339_n, n3339, n3340_n, n3340, n3341_n, n3341, n3342_n, n3342, n3343_n, n3343, n3344_n, n3344, n3345_n, n3345, n3346_n, n3346, n3347_n, n3347, n3348_n, n3348,
 n3349_n, n3349, n3350_n, n3350, n3351_n, n3351, n3352_n, n3352, n3353_n, n3353, n3354_n, n3354, n3355_n, n3355, n3356_n, n3356, n3357_n, n3357, n3358_n, n3358,
 n3359_n, n3359, n3360_n, n3360, n3361_n, n3361, n3362_n, n3362, n3363_n, n3363, n3364_n, n3364, n3365_n, n3365, n3366_n, n3366, n3367_n, n3367, n3368_n, n3368,
 n3369_n, n3369, n3370_n, n3370, n3371_n, n3371, n3372_n, n3372, n3373_n, n3373, n3374_n, n3374, n3375_n, n3375, n3376_n, n3376, n3377_n, n3377, n3378_n, n3378,
 n3379_n, n3379, n3380_n, n3380, n3381_n, n3381, n3382_n, n3382, n3383_n, n3383, n3384_n, n3384, n3385_n, n3385, n3386_n, n3386, n3387_n, n3387, n3388_n, n3388,
 n3389_n, n3389, n3390_n, n3390, n3391_n, n3391, n3392_n, n3392, n3393_n, n3393, n3394_n, n3394, n3395_n, n3395, n3396_n, n3396, n3397_n, n3397, n3398_n, n3398,
 n3399_n, n3399, n3400_n, n3400, n3401_n, n3401, n3402_n, n3402, n3403_n, n3403, n3404_n, n3404, n3405_n, n3405, n3406_n, n3406, n3407_n, n3407, n3408_n, n3408,
 n3409_n, n3409, n3410_n, n3410, n3411_n, n3411, n3412_n, n3412, n3413_n, n3413, n3414_n, n3414, n3415_n, n3415, n3416_n, n3416, n3417_n, n3417, n3418_n, n3418,
 n3419_n, n3419, n3420_n, n3420, n3421_n, n3421, n3422_n, n3422, n3423_n, n3423, n3424_n, n3424, n3425_n, n3425, n3426_n, n3426, n3427_n, n3427, n3428_n, n3428,
 n3429_n, n3429, n3430_n, n3430, n3431_n, n3431, n3432_n, n3432, n3433_n, n3433, n3434_n, n3434, n3435_n, n3435, n3436_n, n3436, n3437_n, n3437, n3438_n, n3438,
 n3439_n, n3439, n3440_n, n3440, n3441_n, n3441, n3442_n, n3442, n3443_n, n3443, n3444_n, n3444, n3445_n, n3445, n3446_n, n3446, n3447_n, n3447, n3448_n, n3448,
 n3449_n, n3449, n3450_n, n3450, n3451_n, n3451, n3452_n, n3452, n3453_n, n3453, n3454_n, n3454, n3455_n, n3455, n3456_n, n3456, n3457_n, n3457, n3458_n, n3458,
 n3459_n;


 wddl_inv U1587 ( .A(n3049), .A_n(n3049_n), .Y_n(n2519_n), .Y(n2519) );
 wddl_inv U1588 ( .A(n2519), .A_n(n2519_n), .Y_n(n2520_n), .Y(n2520) );
 wddl_inv U1589 ( .A(n2995), .A_n(n2995_n), .Y_n(n2521_n), .Y(n2521) );
 wddl_inv U1590 ( .A(n2521), .A_n(n2521_n), .Y_n(n2522_n), .Y(n2522) );
 wddl_inv U1591 ( .A(n3250), .A_n(n3250_n), .Y_n(n2523_n), .Y(n2523) );
 wddl_inv U1592 ( .A(n2523), .A_n(n2523_n), .Y_n(n2524_n), .Y(n2524) );
 wddl_inv U1593 ( .A(n2897), .A_n(n2897_n), .Y_n(n2525_n), .Y(n2525) );
 wddl_inv U1594 ( .A(n2525), .A_n(n2525_n), .Y_n(n2526_n), .Y(n2526) );
 wddl_inv U1595 ( .A(n3299), .A_n(n3299_n), .Y_n(n2527_n), .Y(n2527) );
 wddl_inv U1596 ( .A(n2527), .A_n(n2527_n), .Y_n(n2528_n), .Y(n2528) );
 wddl_inv U1597 ( .A(n2875), .A_n(n2875_n), .Y_n(n2529_n), .Y(n2529) );
 wddl_inv U1598 ( .A(n2529), .A_n(n2529_n), .Y_n(n2530_n), .Y(n2530) );
 wddl_inv U1599 ( .A(n3380), .A_n(n3380_n), .Y_n(n2531_n), .Y(n2531) );
 wddl_inv U1600 ( .A(n2758), .A_n(n2758_n), .Y_n(n2532_n), .Y(n2532) );
 wddl_inv U1601 ( .A(n2532), .A_n(n2532_n), .Y_n(n2533_n), .Y(n2533) );
 wddl_inv U1602 ( .A(n3424), .A_n(n3424_n), .Y_n(n2534_n), .Y(n2534) );
 wddl_inv U1603 ( .A(n2700), .A_n(n2700_n), .Y_n(n2535_n), .Y(n2535) );
 wddl_inv U1604 ( .A(n2535), .A_n(n2535_n), .Y_n(n2536_n), .Y(n2536) );
 wddl_inv U1605 ( .A(n2695), .A_n(n2695_n), .Y_n(n2537_n), .Y(n2537) );
 wddl_inv U1606 ( .A(n2537), .A_n(n2537_n), .Y_n(n2538_n), .Y(n2538) );
 wddl_inv U1607 ( .A(n2690), .A_n(n2690_n), .Y_n(n2539_n), .Y(n2539) );
 wddl_inv U1608 ( .A(n2539), .A_n(n2539_n), .Y_n(n2540_n), .Y(n2540) );
 wddl_inv U1609 ( .A(n2685), .A_n(n2685_n), .Y_n(n2541_n), .Y(n2541) );
 wddl_inv U1610 ( .A(n2541), .A_n(n2541_n), .Y_n(n2542_n), .Y(n2542) );
 wddl_inv U1611 ( .A(n2680), .A_n(n2680_n), .Y_n(n2543_n), .Y(n2543) );
 wddl_inv U1612 ( .A(n2543), .A_n(n2543_n), .Y_n(n2544_n), .Y(n2544) );
 wddl_inv U1613 ( .A(n2676), .A_n(n2676_n), .Y_n(n2545_n), .Y(n2545) );
 wddl_inv U1614 ( .A(n2545), .A_n(n2545_n), .Y_n(n2546_n), .Y(n2546) );
 wddl_inv U1615 ( .A(n2670), .A_n(n2670_n), .Y_n(n2547_n), .Y(n2547) );
 wddl_inv U1616 ( .A(n2547), .A_n(n2547_n), .Y_n(n2548_n), .Y(n2548) );
 wddl_inv U1617 ( .A(n2665), .A_n(n2665_n), .Y_n(n2549_n), .Y(n2549) );
 wddl_inv U1618 ( .A(n2549), .A_n(n2549_n), .Y_n(n2550_n), .Y(n2550) );
 wddl_inv U1619 ( .A(n2710), .A_n(n2710_n), .Y_n(n2551_n), .Y(n2551) );
 wddl_inv U1620 ( .A(n2551), .A_n(n2551_n), .Y_n(n2552_n), .Y(n2552) );
 wddl_inv U1621 ( .A(n2704), .A_n(n2704_n), .Y_n(n2553_n), .Y(n2553) );
 wddl_inv U1622 ( .A(n2553), .A_n(n2553_n), .Y_n(n2554_n), .Y(n2554) );
 wddl_inv U1623 ( .A(n2553), .A_n(n2553_n), .Y_n(n2555_n), .Y(n2555) );
 wddl_inv U1624 ( .A(n2746), .A_n(n2746_n), .Y_n(n2556_n), .Y(n2556) );
 wddl_inv U1625 ( .A(n2556), .A_n(n2556_n), .Y_n(n2557_n), .Y(n2557) );
 wddl_inv U1626 ( .A(n2556), .A_n(n2556_n), .Y_n(n2558_n), .Y(n2558) );
 wddl_inv U1627 ( .A(n2556), .A_n(n2556_n), .Y_n(n2559_n), .Y(n2559) );
 wddl_inv U1628 ( .A(n2835), .A_n(n2835_n), .Y_n(n2560_n), .Y(n2560) );
 wddl_inv U1629 ( .A(n2560), .A_n(n2560_n), .Y_n(n2561_n), .Y(n2561) );
 wddl_inv U1630 ( .A(n2560), .A_n(n2560_n), .Y_n(n2562_n), .Y(n2562) );
 wddl_inv U1631 ( .A(n2560), .A_n(n2560_n), .Y_n(n2563_n), .Y(n2563) );
 wddl_inv U1632 ( .A(n2759), .A_n(n2759_n), .Y_n(n2564_n), .Y(n2564) );
 wddl_inv U1633 ( .A(n2564), .A_n(n2564_n), .Y_n(n2565_n), .Y(n2565) );
 wddl_inv U1634 ( .A(n2564), .A_n(n2564_n), .Y_n(n2566_n), .Y(n2566) );
 wddl_inv U1635 ( .A(n2564), .A_n(n2564_n), .Y_n(n2567_n), .Y(n2567) );
 wddl_inv U1636 ( .A(n2796), .A_n(n2796_n), .Y_n(n2568_n), .Y(n2568) );
 wddl_inv U1637 ( .A(n2568), .A_n(n2568_n), .Y_n(n2569_n), .Y(n2569) );
 wddl_inv U1638 ( .A(n2568), .A_n(n2568_n), .Y_n(n2570_n), .Y(n2570) );
 wddl_inv U1639 ( .A(n2568), .A_n(n2568_n), .Y_n(n2571_n), .Y(n2571) );
 wddl_inv U1640 ( .A(n2762), .A_n(n2762_n), .Y_n(n2572_n), .Y(n2572) );
 wddl_inv U1641 ( .A(n2572), .A_n(n2572_n), .Y_n(n2573_n), .Y(n2573) );
 wddl_inv U1642 ( .A(n2572), .A_n(n2572_n), .Y_n(n2576_n), .Y(n2576) );
 wddl_inv U1643 ( .A(n2572), .A_n(n2572_n), .Y_n(n2574_n), .Y(n2574) );
 wddl_inv U1644 ( .A(n2572), .A_n(n2572_n), .Y_n(n2575_n), .Y(n2575) );
 wddl_inv U1645 ( .A(n2798), .A_n(n2798_n), .Y_n(n2577_n), .Y(n2577) );
 wddl_inv U1646 ( .A(n2577), .A_n(n2577_n), .Y_n(n2578_n), .Y(n2578) );
 wddl_inv U1647 ( .A(n2577), .A_n(n2577_n), .Y_n(n2581_n), .Y(n2581) );
 wddl_inv U1648 ( .A(n2577), .A_n(n2577_n), .Y_n(n2579_n), .Y(n2579) );
 wddl_inv U1649 ( .A(n2577), .A_n(n2577_n), .Y_n(n2580_n), .Y(n2580) );
 wddl_inv U1650 ( .A(n2757), .A_n(n2757_n), .Y_n(n2582_n), .Y(n2582) );
 wddl_inv U1651 ( .A(n2582), .A_n(n2582_n), .Y_n(n2583_n), .Y(n2583) );
 wddl_inv U1652 ( .A(n2582), .A_n(n2582_n), .Y_n(n2586_n), .Y(n2586) );
 wddl_inv U1653 ( .A(n2582), .A_n(n2582_n), .Y_n(n2584_n), .Y(n2584) );
 wddl_inv U1654 ( .A(n2582), .A_n(n2582_n), .Y_n(n2585_n), .Y(n2585) );
 wddl_inv U1655 ( .A(n2868), .A_n(n2868_n), .Y_n(n2587_n), .Y(n2587) );
 wddl_inv U1656 ( .A(n2587), .A_n(n2587_n), .Y_n(n2588_n), .Y(n2588) );
 wddl_inv U1657 ( .A(n2587), .A_n(n2587_n), .Y_n(n2591_n), .Y(n2591) );
 wddl_inv U1658 ( .A(n2587), .A_n(n2587_n), .Y_n(n2589_n), .Y(n2589) );
 wddl_inv U1659 ( .A(n2587), .A_n(n2587_n), .Y_n(n2590_n), .Y(n2590) );
 wddl_inv U1660 ( .A(n2743), .A_n(n2743_n), .Y_n(n2592_n), .Y(n2592) );
 wddl_inv U1661 ( .A(n2592), .A_n(n2592_n), .Y_n(n2593_n), .Y(n2593) );
 wddl_inv U1662 ( .A(n2592), .A_n(n2592_n), .Y_n(n2596_n), .Y(n2596) );
 wddl_inv U1663 ( .A(n2592), .A_n(n2592_n), .Y_n(n2594_n), .Y(n2594) );
 wddl_inv U1664 ( .A(n2592), .A_n(n2592_n), .Y_n(n2595_n), .Y(n2595) );
 wddl_inv U1665 ( .A(n2822), .A_n(n2822_n), .Y_n(n2597_n), .Y(n2597) );
 wddl_inv U1666 ( .A(n2597), .A_n(n2597_n), .Y_n(n2598_n), .Y(n2598) );
 wddl_inv U1667 ( .A(n2597), .A_n(n2597_n), .Y_n(n2601_n), .Y(n2601) );
 wddl_inv U1668 ( .A(n2597), .A_n(n2597_n), .Y_n(n2599_n), .Y(n2599) );
 wddl_inv U1669 ( .A(n2597), .A_n(n2597_n), .Y_n(n2600_n), .Y(n2600) );
 wddl_inv U1670 ( .A(n2771), .A_n(n2771_n), .Y_n(n2602_n), .Y(n2602) );
 wddl_inv U1671 ( .A(n2602), .A_n(n2602_n), .Y_n(n2603_n), .Y(n2603) );
 wddl_inv U1672 ( .A(n2602), .A_n(n2602_n), .Y_n(n2606_n), .Y(n2606) );
 wddl_inv U1673 ( .A(n2602), .A_n(n2602_n), .Y_n(n2604_n), .Y(n2604) );
 wddl_inv U1674 ( .A(n2602), .A_n(n2602_n), .Y_n(n2605_n), .Y(n2605) );
 wddl_inv U1675 ( .A(n2829), .A_n(n2829_n), .Y_n(n2607_n), .Y(n2607) );
 wddl_inv U1676 ( .A(n2607), .A_n(n2607_n), .Y_n(n2608_n), .Y(n2608) );
 wddl_inv U1677 ( .A(n2607), .A_n(n2607_n), .Y_n(n2611_n), .Y(n2611) );
 wddl_inv U1678 ( .A(n2607), .A_n(n2607_n), .Y_n(n2609_n), .Y(n2609) );
 wddl_inv U1679 ( .A(n2607), .A_n(n2607_n), .Y_n(n2610_n), .Y(n2610) );
 wddl_inv U1680 ( .A(n2748), .A_n(n2748_n), .Y_n(n2612_n), .Y(n2612) );
 wddl_inv U1681 ( .A(n2612), .A_n(n2612_n), .Y_n(n2613_n), .Y(n2613) );
 wddl_inv U1682 ( .A(n2612), .A_n(n2612_n), .Y_n(n2616_n), .Y(n2616) );
 wddl_inv U1683 ( .A(n2612), .A_n(n2612_n), .Y_n(n2614_n), .Y(n2614) );
 wddl_inv U1684 ( .A(n2612), .A_n(n2612_n), .Y_n(n2615_n), .Y(n2615) );
 wddl_inv U1685 ( .A(n2874), .A_n(n2874_n), .Y_n(n2617_n), .Y(n2617) );
 wddl_inv U1686 ( .A(n2617), .A_n(n2617_n), .Y_n(n2618_n), .Y(n2618) );
 wddl_inv U1687 ( .A(n2617), .A_n(n2617_n), .Y_n(n2621_n), .Y(n2621) );
 wddl_inv U1688 ( .A(n2617), .A_n(n2617_n), .Y_n(n2619_n), .Y(n2619) );
 wddl_inv U1689 ( .A(n2617), .A_n(n2617_n), .Y_n(n2620_n), .Y(n2620) );
 wddl_inv U1690 ( .A(n2770), .A_n(n2770_n), .Y_n(n2622_n), .Y(n2622) );
 wddl_inv U1691 ( .A(n2622), .A_n(n2622_n), .Y_n(n2623_n), .Y(n2623) );
 wddl_inv U1692 ( .A(n2622), .A_n(n2622_n), .Y_n(n2626_n), .Y(n2626) );
 wddl_inv U1693 ( .A(n2622), .A_n(n2622_n), .Y_n(n2624_n), .Y(n2624) );
 wddl_inv U1694 ( .A(n2622), .A_n(n2622_n), .Y_n(n2625_n), .Y(n2625) );
 wddl_inv U1695 ( .A(n2773), .A_n(n2773_n), .Y_n(n2627_n), .Y(n2627) );
 wddl_inv U1696 ( .A(n2627), .A_n(n2627_n), .Y_n(n2628_n), .Y(n2628) );
 wddl_inv U1697 ( .A(n2627), .A_n(n2627_n), .Y_n(n2631_n), .Y(n2631) );
 wddl_inv U1698 ( .A(n2627), .A_n(n2627_n), .Y_n(n2629_n), .Y(n2629) );
 wddl_inv U1699 ( .A(n2627), .A_n(n2627_n), .Y_n(n2630_n), .Y(n2630) );
 wddl_inv U1700 ( .A(n2764), .A_n(n2764_n), .Y_n(n2632_n), .Y(n2632) );
 wddl_inv U1701 ( .A(n2632), .A_n(n2632_n), .Y_n(n2633_n), .Y(n2633) );
 wddl_inv U1702 ( .A(n2632), .A_n(n2632_n), .Y_n(n2636_n), .Y(n2636) );
 wddl_inv U1703 ( .A(n2632), .A_n(n2632_n), .Y_n(n2634_n), .Y(n2634) );
 wddl_inv U1704 ( .A(n2632), .A_n(n2632_n), .Y_n(n2635_n), .Y(n2635) );
 wddl_inv U1705 ( .A(n2797), .A_n(n2797_n), .Y_n(n2637_n), .Y(n2637) );
 wddl_inv U1706 ( .A(n2637), .A_n(n2637_n), .Y_n(n2638_n), .Y(n2638) );
 wddl_inv U1707 ( .A(n2637), .A_n(n2637_n), .Y_n(n2641_n), .Y(n2641) );
 wddl_inv U1708 ( .A(n2637), .A_n(n2637_n), .Y_n(n2639_n), .Y(n2639) );
 wddl_inv U1709 ( .A(n2637), .A_n(n2637_n), .Y_n(n2640_n), .Y(n2640) );
 wddl_inv U1710 ( .A(n2741), .A_n(n2741_n), .Y_n(n2642_n), .Y(n2642) );
 wddl_inv U1711 ( .A(n2642), .A_n(n2642_n), .Y_n(n2643_n), .Y(n2643) );
 wddl_inv U1712 ( .A(n2642), .A_n(n2642_n), .Y_n(n2646_n), .Y(n2646) );
 wddl_inv U1713 ( .A(n2642), .A_n(n2642_n), .Y_n(n2644_n), .Y(n2644) );
 wddl_inv U1714 ( .A(n2642), .A_n(n2642_n), .Y_n(n2645_n), .Y(n2645) );
 wddl_inv U1715 ( .A(n2760), .A_n(n2760_n), .Y_n(n2647_n), .Y(n2647) );
 wddl_inv U1716 ( .A(n2647), .A_n(n2647_n), .Y_n(n2648_n), .Y(n2648) );
 wddl_inv U1717 ( .A(n2647), .A_n(n2647_n), .Y_n(n2651_n), .Y(n2651) );
 wddl_inv U1718 ( .A(n2647), .A_n(n2647_n), .Y_n(n2649_n), .Y(n2649) );
 wddl_inv U1719 ( .A(n2647), .A_n(n2647_n), .Y_n(n2650_n), .Y(n2650) );
 wddl_inv U1720 ( .A(n2749), .A_n(n2749_n), .Y_n(n2652_n), .Y(n2652) );
 wddl_inv U1721 ( .A(n2652), .A_n(n2652_n), .Y_n(n2653_n), .Y(n2653) );
 wddl_inv U1722 ( .A(n2652), .A_n(n2652_n), .Y_n(n2656_n), .Y(n2656) );
 wddl_inv U1723 ( .A(n2652), .A_n(n2652_n), .Y_n(n2654_n), .Y(n2654) );
 wddl_inv U1724 ( .A(n2652), .A_n(n2652_n), .Y_n(n2655_n), .Y(n2655) );
 wddl_inv U1725 ( .A(n2811), .A_n(n2811_n), .Y_n(n2657_n), .Y(n2657) );
 wddl_inv U1726 ( .A(n2657), .A_n(n2657_n), .Y_n(n2658_n), .Y(n2658) );
 wddl_inv U1727 ( .A(n2657), .A_n(n2657_n), .Y_n(n2661_n), .Y(n2661) );
 wddl_inv U1728 ( .A(n2657), .A_n(n2657_n), .Y_n(n2659_n), .Y(n2659) );
 wddl_inv U1729 ( .A(n2657), .A_n(n2657_n), .Y_n(n2660_n), .Y(n2660) );
 wddl_inv U1730 ( .A(n2786), .A_n(n2786_n), .Y_n(n2662_n), .Y(n2662) );
 wddl_inv U1731 ( .A(n2662), .A_n(n2662_n), .Y_n(n2663_n), .Y(n2663) );
 wddl_inv U1732 ( .A(n2662), .A_n(n2662_n), .Y_n(n2666_n), .Y(n2666) );
 wddl_inv U1733 ( .A(n2662), .A_n(n2662_n), .Y_n(n2664_n), .Y(n2664) );
 wddl_inv U1734 ( .A(n2662), .A_n(n2662_n), .Y_n(n2665_n), .Y(n2665) );
 wddl_inv U1735 ( .A(n2788), .A_n(n2788_n), .Y_n(n2667_n), .Y(n2667) );
 wddl_inv U1736 ( .A(n2667), .A_n(n2667_n), .Y_n(n2668_n), .Y(n2668) );
 wddl_inv U1737 ( .A(n2667), .A_n(n2667_n), .Y_n(n2671_n), .Y(n2671) );
 wddl_inv U1738 ( .A(n2667), .A_n(n2667_n), .Y_n(n2669_n), .Y(n2669) );
 wddl_inv U1739 ( .A(n2667), .A_n(n2667_n), .Y_n(n2670_n), .Y(n2670) );
 wddl_inv U1740 ( .A(n2772), .A_n(n2772_n), .Y_n(n2672_n), .Y(n2672) );
 wddl_inv U1741 ( .A(n2672), .A_n(n2672_n), .Y_n(n2673_n), .Y(n2673) );
 wddl_inv U1742 ( .A(n2672), .A_n(n2672_n), .Y_n(n2676_n), .Y(n2676) );
 wddl_inv U1743 ( .A(n2672), .A_n(n2672_n), .Y_n(n2674_n), .Y(n2674) );
 wddl_inv U1744 ( .A(n2672), .A_n(n2672_n), .Y_n(n2675_n), .Y(n2675) );
 wddl_inv U1745 ( .A(n2804), .A_n(n2804_n), .Y_n(n2677_n), .Y(n2677) );
 wddl_inv U1746 ( .A(n2677), .A_n(n2677_n), .Y_n(n2678_n), .Y(n2678) );
 wddl_inv U1747 ( .A(n2677), .A_n(n2677_n), .Y_n(n2681_n), .Y(n2681) );
 wddl_inv U1748 ( .A(n2677), .A_n(n2677_n), .Y_n(n2679_n), .Y(n2679) );
 wddl_inv U1749 ( .A(n2677), .A_n(n2677_n), .Y_n(n2680_n), .Y(n2680) );
 wddl_inv U1750 ( .A(n2756), .A_n(n2756_n), .Y_n(n2682_n), .Y(n2682) );
 wddl_inv U1751 ( .A(n2682), .A_n(n2682_n), .Y_n(n2683_n), .Y(n2683) );
 wddl_inv U1752 ( .A(n2682), .A_n(n2682_n), .Y_n(n2686_n), .Y(n2686) );
 wddl_inv U1753 ( .A(n2682), .A_n(n2682_n), .Y_n(n2684_n), .Y(n2684) );
 wddl_inv U1754 ( .A(n2682), .A_n(n2682_n), .Y_n(n2685_n), .Y(n2685) );
 wddl_inv U1755 ( .A(n2830), .A_n(n2830_n), .Y_n(n2687_n), .Y(n2687) );
 wddl_inv U1756 ( .A(n2687), .A_n(n2687_n), .Y_n(n2688_n), .Y(n2688) );
 wddl_inv U1757 ( .A(n2687), .A_n(n2687_n), .Y_n(n2691_n), .Y(n2691) );
 wddl_inv U1758 ( .A(n2687), .A_n(n2687_n), .Y_n(n2689_n), .Y(n2689) );
 wddl_inv U1759 ( .A(n2687), .A_n(n2687_n), .Y_n(n2690_n), .Y(n2690) );
 wddl_inv U1760 ( .A(n2744), .A_n(n2744_n), .Y_n(n2692_n), .Y(n2692) );
 wddl_inv U1761 ( .A(n2692), .A_n(n2692_n), .Y_n(n2693_n), .Y(n2693) );
 wddl_inv U1762 ( .A(n2692), .A_n(n2692_n), .Y_n(n2696_n), .Y(n2696) );
 wddl_inv U1763 ( .A(n2692), .A_n(n2692_n), .Y_n(n2694_n), .Y(n2694) );
 wddl_inv U1764 ( .A(n2692), .A_n(n2692_n), .Y_n(n2695_n), .Y(n2695) );
 wddl_inv U1765 ( .A(n2895), .A_n(n2895_n), .Y_n(n2697_n), .Y(n2697) );
 wddl_inv U1766 ( .A(n2697), .A_n(n2697_n), .Y_n(n2698_n), .Y(n2698) );
 wddl_inv U1767 ( .A(n2697), .A_n(n2697_n), .Y_n(n2701_n), .Y(n2701) );
 wddl_inv U1768 ( .A(n2697), .A_n(n2697_n), .Y_n(n2699_n), .Y(n2699) );
 wddl_inv U1769 ( .A(n2697), .A_n(n2697_n), .Y_n(n2700_n), .Y(n2700) );
 wddl_inv U1770 ( .A(n2805), .A_n(n2805_n), .Y_n(n2702_n), .Y(n2702) );
 wddl_inv U1771 ( .A(n2702), .A_n(n2702_n), .Y_n(n2703_n), .Y(n2703) );
 wddl_inv U1772 ( .A(n2702), .A_n(n2702_n), .Y_n(n2705_n), .Y(n2705) );
 wddl_inv U1773 ( .A(n2702), .A_n(n2702_n), .Y_n(n2704_n), .Y(n2704) );
 wddl_inv U1774 ( .A(n2799), .A_n(n2799_n), .Y_n(n2706_n), .Y(n2706) );
 wddl_inv U1775 ( .A(n2706), .A_n(n2706_n), .Y_n(n2707_n), .Y(n2707) );
 wddl_inv U1776 ( .A(n2706), .A_n(n2706_n), .Y_n(n2710_n), .Y(n2710) );
 wddl_inv U1777 ( .A(n2706), .A_n(n2706_n), .Y_n(n2708_n), .Y(n2708) );
 wddl_inv U1778 ( .A(n2706), .A_n(n2706_n), .Y_n(n2709_n), .Y(n2709) );
 wddl_inv U1779 ( .A(a[4]), .A_n(a_n[4]), .Y_n(n2711_n), .Y(n2711) );
 wddl_inv U1780 ( .A(n2711), .A_n(n2711_n), .Y_n(n2712_n), .Y(n2712) );
 wddl_inv U1781 ( .A(a[6]), .A_n(a_n[6]), .Y_n(n2713_n), .Y(n2713) );
 wddl_inv U1782 ( .A(n2713), .A_n(n2713_n), .Y_n(n2714_n), .Y(n2714) );
 wddl_inv U1783 ( .A(a[2]), .A_n(a_n[2]), .Y_n(n2715_n), .Y(n2715) );
 wddl_inv U1784 ( .A(n2715), .A_n(n2715_n), .Y_n(n2716_n), .Y(n2716) );
 wddl_inv U1785 ( .A(a[1]), .A_n(a_n[1]), .Y_n(n2717_n), .Y(n2717) );
 wddl_inv U1786 ( .A(n2717), .A_n(n2717_n), .Y_n(n2718_n), .Y(n2718) );
 wddl_inv U1787 ( .A(a[3]), .A_n(a_n[3]), .Y_n(n2719_n), .Y(n2719) );
 wddl_inv U1788 ( .A(n2719), .A_n(n2719_n), .Y_n(n2720_n), .Y(n2720) );
 wddl_inv U1789 ( .A(a[7]), .A_n(a_n[7]), .Y_n(n2721_n), .Y(n2721) );
 wddl_inv U1790 ( .A(n2721), .A_n(n2721_n), .Y_n(n2722_n), .Y(n2722) );
 wddl_inv U1791 ( .A(a[5]), .A_n(a_n[5]), .Y_n(n2723_n), .Y(n2723) );
 wddl_inv U1792 ( .A(n2723), .A_n(n2723_n), .Y_n(n2724_n), .Y(n2724) );
 wddl_inv U1793 ( .A(a[0]), .A_n(a_n[0]), .Y_n(n2725_n), .Y(n2725) );
 wddl_inv U1794 ( .A(n2725), .A_n(n2725_n), .Y_n(n2726_n), .Y(n2726) );
 wddl_or U1795 ( .A(n3028), .A_n(n3028_n), .B(n3285), .B_n(n3285_n), .Y_n(d_n[0]), .Y(d[0]) );
 wddl_or U1796 ( .A(n3286), .A_n(n3286_n), .B(n3287), .B_n(n3287_n), .Y_n(n3285_n), .Y(n3285) );
 wddl_or U1797 ( .A(n3004), .A_n(n3004_n), .B(n3288), .B_n(n3288_n), .Y_n(n3287_n), .Y(n3287) );
 wddl_or U1798 ( .A(n3289), .A_n(n3289_n), .B(n3290), .B_n(n3290_n), .Y_n(n3288_n), .Y(n3288) );
 wddl_or U1799 ( .A(n3291), .A_n(n3291_n), .B(n3292), .B_n(n3292_n), .Y_n(n3290_n), .Y(n3290) );
 wddl_or U1800 ( .A(n3293), .A_n(n3293_n), .B(n3294), .B_n(n3294_n), .Y_n(n3292_n), .Y(n3292) );
 wddl_and U1801 ( .A(n2773), .A_n(n2773_n), .B(n2664), .B_n(n2664_n), .Y_n(n3294_n), .Y(n3294) );
 wddl_and U1802 ( .A(n2614), .A_n(n2614_n), .B(n2789), .B_n(n2789_n), .Y_n(n3293_n), .Y(n3293) );
 wddl_or U1803 ( .A(n3295), .A_n(n3295_n), .B(n3296), .B_n(n3296_n), .Y_n(n3291_n), .Y(n3291) );
 wddl_and U1804 ( .A(n2569), .A_n(n2569_n), .B(n3297), .B_n(n3297_n), .Y_n(n3296_n), .Y(n3296) );
 wddl_or U1805 ( .A(n2554), .A_n(n2554_n), .B(n2526), .B_n(n2526_n), .Y_n(n3297_n), .Y(n3297) );
 wddl_and U1806 ( .A(n2598), .A_n(n2598_n), .B(n3298), .B_n(n3298_n), .Y_n(n3295_n), .Y(n3295) );
 wddl_and U1807 ( .A(n2714), .A_n(n2714_n), .B(n2528), .B_n(n2528_n), .Y_n(n3298_n), .Y(n3298) );
 wddl_or U1808 ( .A(n3300), .A_n(n3300_n), .B(n3301), .B_n(n3301_n), .Y_n(n3289_n), .Y(n3289) );
 wddl_or U1809 ( .A(n2884), .A_n(n2884_n), .B(n3302), .B_n(n3302_n), .Y_n(n3301_n), .Y(n3301) );
 wddl_or U1810 ( .A(n3303), .A_n(n3303_n), .B(n3304), .B_n(n3304_n), .Y_n(n3302_n), .Y(n3302) );
 wddl_or U1811 ( .A(n3305), .A_n(n3305_n), .B(n3306), .B_n(n3306_n), .Y_n(n3304_n), .Y(n3304) );
 wddl_and U1812 ( .A(n2685), .A_n(n2685_n), .B(n2764), .B_n(n2764_n), .Y_n(n3305_n), .Y(n3305) );
 wddl_and U1813 ( .A(n2604), .A_n(n2604_n), .B(n2869), .B_n(n2869_n), .Y_n(n3303_n), .Y(n3303) );
 wddl_or U1814 ( .A(n2828), .A_n(n2828_n), .B(n3307), .B_n(n3307_n), .Y_n(n3300_n), .Y(n3300) );
 wddl_and U1815 ( .A(n2562), .A_n(n2562_n), .B(n2520), .B_n(n2520_n), .Y_n(n3307_n), .Y(n3307) );
 wddl_or U1816 ( .A(n2870), .A_n(n2870_n), .B(n2983), .B_n(n2983_n), .Y_n(n3286_n), .Y(n3286) );
 wddl_or U1817 ( .A(n2727), .A_n(n2727_n), .B(n2774), .B_n(n2774_n), .Y_n(d_n[6]), .Y(d[6]) );
 wddl_or U1818 ( .A(n2775), .A_n(n2775_n), .B(n2776), .B_n(n2776_n), .Y_n(n2774_n), .Y(n2774) );
 wddl_or U1819 ( .A(n2777), .A_n(n2777_n), .B(n2778), .B_n(n2778_n), .Y_n(n2776_n), .Y(n2776) );
 wddl_or U1820 ( .A(n2779), .A_n(n2779_n), .B(n2780), .B_n(n2780_n), .Y_n(n2778_n), .Y(n2778) );
 wddl_or U1821 ( .A(n2781), .A_n(n2781_n), .B(n2782), .B_n(n2782_n), .Y_n(n2780_n), .Y(n2780) );
 wddl_or U1822 ( .A(n2783), .A_n(n2783_n), .B(n2784), .B_n(n2784_n), .Y_n(n2782_n), .Y(n2782) );
 wddl_and U1823 ( .A(n2673), .A_n(n2673_n), .B(n2785), .B_n(n2785_n), .Y_n(n2784_n), .Y(n2784) );
 wddl_and U1824 ( .A(n2666), .A_n(n2666_n), .B(n2787), .B_n(n2787_n), .Y_n(n2783_n), .Y(n2783) );
 wddl_or U1825 ( .A(n2548), .A_n(n2548_n), .B(n2789), .B_n(n2789_n), .Y_n(n2787_n), .Y(n2787) );
 wddl_or U1826 ( .A(n2591), .A_n(n2591_n), .B(n2557), .B_n(n2557_n), .Y_n(n2789_n), .Y(n2789) );
 wddl_or U1827 ( .A(n2790), .A_n(n2790_n), .B(n2791), .B_n(n2791_n), .Y_n(n2781_n), .Y(n2781) );
 wddl_or U1828 ( .A(n2792), .A_n(n2792_n), .B(n2793), .B_n(n2793_n), .Y_n(n2791_n), .Y(n2791) );
 wddl_or U1829 ( .A(n2794), .A_n(n2794_n), .B(n2795), .B_n(n2795_n), .Y_n(n2793_n), .Y(n2793) );
 wddl_and U1830 ( .A(n2571), .A_n(n2571_n), .B(n2640), .B_n(n2640_n), .Y_n(n2795_n), .Y(n2795) );
 wddl_and U1831 ( .A(n2579), .A_n(n2579_n), .B(n2585), .B_n(n2585_n), .Y_n(n2794_n), .Y(n2794) );
 wddl_and U1832 ( .A(n2552), .A_n(n2552_n), .B(n2800), .B_n(n2800_n), .Y_n(n2792_n), .Y(n2792) );
 wddl_or U1833 ( .A(n2801), .A_n(n2801_n), .B(n2802), .B_n(n2802_n), .Y_n(n2790_n), .Y(n2790) );
 wddl_and U1834 ( .A(n2625), .A_n(n2625_n), .B(n2803), .B_n(n2803_n), .Y_n(n2802_n), .Y(n2802) );
 wddl_or U1835 ( .A(n2684), .A_n(n2684_n), .B(n2681), .B_n(n2681_n), .Y_n(n2803_n), .Y(n2803) );
 wddl_and U1836 ( .A(n2704), .A_n(n2704_n), .B(n2806), .B_n(n2806_n), .Y_n(n2801_n), .Y(n2801) );
 wddl_or U1837 ( .A(n2633), .A_n(n2633_n), .B(n2538), .B_n(n2538_n), .Y_n(n2806_n), .Y(n2806) );
 wddl_or U1838 ( .A(n2807), .A_n(n2807_n), .B(n2808), .B_n(n2808_n), .Y_n(n2775_n), .Y(n2775) );
 wddl_or U1839 ( .A(n2809), .A_n(n2809_n), .B(n2810), .B_n(n2810_n), .Y_n(n2808_n), .Y(n2808) );
 wddl_and U1840 ( .A(n2771), .A_n(n2771_n), .B(n2659), .B_n(n2659_n), .Y_n(n2810_n), .Y(n2810) );
 wddl_or U1841 ( .A(n2844), .A_n(n2844_n), .B(n2845), .B_n(n2845_n), .Y_n(d_n[5]), .Y(d[5]) );
 wddl_or U1842 ( .A(n2846), .A_n(n2846_n), .B(n2847), .B_n(n2847_n), .Y_n(n2845_n), .Y(n2845) );
 wddl_or U1843 ( .A(n2848), .A_n(n2848_n), .B(n2849), .B_n(n2849_n), .Y_n(n2847_n), .Y(n2847) );
 wddl_or U1844 ( .A(n2850), .A_n(n2850_n), .B(n2851), .B_n(n2851_n), .Y_n(n2849_n), .Y(n2849) );
 wddl_or U1845 ( .A(n2852), .A_n(n2852_n), .B(n2853), .B_n(n2853_n), .Y_n(n2850_n), .Y(n2850) );
 wddl_or U1846 ( .A(n2854), .A_n(n2854_n), .B(n2855), .B_n(n2855_n), .Y_n(n2853_n), .Y(n2853) );
 wddl_and U1847 ( .A(n2566), .A_n(n2566_n), .B(n2856), .B_n(n2856_n), .Y_n(n2855_n), .Y(n2855) );
 wddl_and U1848 ( .A(n2835), .A_n(n2835_n), .B(n2857), .B_n(n2857_n), .Y_n(n2854_n), .Y(n2854) );
 wddl_or U1849 ( .A(n2624), .A_n(n2624_n), .B(n2695), .B_n(n2695_n), .Y_n(n2857_n), .Y(n2857) );
 wddl_or U1850 ( .A(n2858), .A_n(n2858_n), .B(n2859), .B_n(n2859_n), .Y_n(n2852_n), .Y(n2852) );
 wddl_or U1851 ( .A(n2860), .A_n(n2860_n), .B(n2861), .B_n(n2861_n), .Y_n(n2859_n), .Y(n2859) );
 wddl_and U1852 ( .A(n2656), .A_n(n2656_n), .B(n2862), .B_n(n2862_n), .Y_n(n2861_n), .Y(n2861) );
 wddl_and U1853 ( .A(n2786), .A_n(n2786_n), .B(n2785), .B_n(n2785_n), .Y_n(n2860_n), .Y(n2860) );
 wddl_or U1854 ( .A(n2605), .A_n(n2605_n), .B(n2863), .B_n(n2863_n), .Y_n(n2785_n), .Y(n2785) );
 wddl_or U1855 ( .A(n2864), .A_n(n2864_n), .B(n2865), .B_n(n2865_n), .Y_n(n2858_n), .Y(n2858) );
 wddl_or U1856 ( .A(n2866), .A_n(n2866_n), .B(n2867), .B_n(n2867_n), .Y_n(n2865_n), .Y(n2865) );
 wddl_and U1857 ( .A(n2542), .A_n(n2542_n), .B(n2760), .B_n(n2760_n), .Y_n(n2867_n), .Y(n2867) );
 wddl_and U1858 ( .A(n2591), .A_n(n2591_n), .B(n2869), .B_n(n2869_n), .Y_n(n2864_n), .Y(n2864) );
 wddl_or U1859 ( .A(n2870), .A_n(n2870_n), .B(n2871), .B_n(n2871_n), .Y_n(n2846_n), .Y(n2846) );
 wddl_or U1860 ( .A(n2872), .A_n(n2872_n), .B(n2873), .B_n(n2873_n), .Y_n(n2871_n), .Y(n2871) );
 wddl_and U1861 ( .A(n2708), .A_n(n2708_n), .B(n2621), .B_n(n2621_n), .Y_n(n2873_n), .Y(n2873) );
 wddl_and U1862 ( .A(n2601), .A_n(n2601_n), .B(n2875), .B_n(n2875_n), .Y_n(n2872_n), .Y(n2872) );
 wddl_or U1863 ( .A(n3344), .A_n(n3344_n), .B(n3345), .B_n(n3345_n), .Y_n(n2870_n), .Y(n2870) );
 wddl_or U1864 ( .A(n3346), .A_n(n3346_n), .B(n3347), .B_n(n3347_n), .Y_n(n3345_n), .Y(n3345) );
 wddl_and U1865 ( .A(n2593), .A_n(n2593_n), .B(n3348), .B_n(n3348_n), .Y_n(n3347_n), .Y(n3347) );
 wddl_or U1866 ( .A(n2704), .A_n(n2704_n), .B(n2691), .B_n(n2691_n), .Y_n(n3348_n), .Y(n3348) );
 wddl_and U1867 ( .A(n2606), .A_n(n2606_n), .B(n3349), .B_n(n3349_n), .Y_n(n3346_n), .Y(n3346) );
 wddl_or U1868 ( .A(n2658), .A_n(n2658_n), .B(n3080), .B_n(n3080_n), .Y_n(n3349_n), .Y(n3349) );
 wddl_or U1869 ( .A(n3350), .A_n(n3350_n), .B(n3351), .B_n(n3351_n), .Y_n(n3344_n), .Y(n3344) );
 wddl_or U1870 ( .A(n3352), .A_n(n3352_n), .B(n3353), .B_n(n3353_n), .Y_n(n3351_n), .Y(n3351) );
 wddl_and U1871 ( .A(n2570), .A_n(n2570_n), .B(n3354), .B_n(n3354_n), .Y_n(n3353_n), .Y(n3353) );
 wddl_or U1872 ( .A(n2756), .A_n(n2756_n), .B(n2576), .B_n(n2576_n), .Y_n(n3354_n), .Y(n3354) );
 wddl_and U1873 ( .A(n2584), .A_n(n2584_n), .B(n3355), .B_n(n3355_n), .Y_n(n3352_n), .Y(n3352) );
 wddl_or U1874 ( .A(n2710), .A_n(n2710_n), .B(n2898), .B_n(n2898_n), .Y_n(n3355_n), .Y(n3355) );
 wddl_or U1875 ( .A(n3356), .A_n(n3356_n), .B(n3357), .B_n(n3357_n), .Y_n(n3350_n), .Y(n3350) );
 wddl_or U1876 ( .A(n3358), .A_n(n3358_n), .B(n3359), .B_n(n3359_n), .Y_n(n3357_n), .Y(n3357) );
 wddl_or U1877 ( .A(n3360), .A_n(n3360_n), .B(n3361), .B_n(n3361_n), .Y_n(n3359_n), .Y(n3359) );
 wddl_and U1878 ( .A(n2579), .A_n(n2579_n), .B(n2744), .B_n(n2744_n), .Y_n(n3361_n), .Y(n3361) );
 wddl_and U1879 ( .A(n2701), .A_n(n2701_n), .B(n2668), .B_n(n2668_n), .Y_n(n3360_n), .Y(n3360) );
 wddl_and U1880 ( .A(n2651), .A_n(n2651_n), .B(n3256), .B_n(n3256_n), .Y_n(n3358_n), .Y(n3358) );
 wddl_and U1881 ( .A(n2618), .A_n(n2618_n), .B(n2912), .B_n(n2912_n), .Y_n(n3356_n), .Y(n3356) );
 wddl_or U1882 ( .A(n2876), .A_n(n2876_n), .B(n2877), .B_n(n2877_n), .Y_n(d_n[4]), .Y(d[4]) );
 wddl_or U1883 ( .A(n2878), .A_n(n2878_n), .B(n2879), .B_n(n2879_n), .Y_n(n2877_n), .Y(n2877) );
 wddl_or U1884 ( .A(n2880), .A_n(n2880_n), .B(n2881), .B_n(n2881_n), .Y_n(n2879_n), .Y(n2879) );
 wddl_or U1885 ( .A(n2882), .A_n(n2882_n), .B(n2883), .B_n(n2883_n), .Y_n(n2881_n), .Y(n2881) );
 wddl_or U1886 ( .A(n2884), .A_n(n2884_n), .B(n2885), .B_n(n2885_n), .Y_n(n2883_n), .Y(n2883) );
 wddl_or U1887 ( .A(n2886), .A_n(n2886_n), .B(n2887), .B_n(n2887_n), .Y_n(n2885_n), .Y(n2885) );
 wddl_and U1888 ( .A(n2563), .A_n(n2563_n), .B(n2749), .B_n(n2749_n), .Y_n(n2887_n), .Y(n2887) );
 wddl_and U1889 ( .A(n2796), .A_n(n2796_n), .B(n2888), .B_n(n2888_n), .Y_n(n2886_n), .Y(n2886) );
 wddl_and U1890 ( .A(n2626), .A_n(n2626_n), .B(n2689), .B_n(n2689_n), .Y_n(n2884_n), .Y(n2884) );
 wddl_or U1891 ( .A(n2889), .A_n(n2889_n), .B(n2890), .B_n(n2890_n), .Y_n(n2882_n), .Y(n2882) );
 wddl_or U1892 ( .A(n2891), .A_n(n2891_n), .B(n2892), .B_n(n2892_n), .Y_n(n2890_n), .Y(n2890) );
 wddl_or U1893 ( .A(n2893), .A_n(n2893_n), .B(n2894), .B_n(n2894_n), .Y_n(n2892_n), .Y(n2892) );
 wddl_and U1894 ( .A(n2704), .A_n(n2704_n), .B(n2786), .B_n(n2786_n), .Y_n(n2894_n), .Y(n2894) );
 wddl_and U1895 ( .A(n2699), .A_n(n2699_n), .B(n2896), .B_n(n2896_n), .Y_n(n2893_n), .Y(n2893) );
 wddl_or U1896 ( .A(n2686), .A_n(n2686_n), .B(n2897), .B_n(n2897_n), .Y_n(n2896_n), .Y(n2896) );
 wddl_and U1897 ( .A(n2659), .A_n(n2659_n), .B(n2898), .B_n(n2898_n), .Y_n(n2891_n), .Y(n2891) );
 wddl_or U1898 ( .A(n2679), .A_n(n2679_n), .B(n2548), .B_n(n2548_n), .Y_n(n2898_n), .Y(n2898) );
 wddl_and U1899 ( .A(n2585), .A_n(n2585_n), .B(n2899), .B_n(n2899_n), .Y_n(n2889_n), .Y(n2889) );
 wddl_or U1900 ( .A(n2671), .A_n(n2671_n), .B(n2900), .B_n(n2900_n), .Y_n(n2899_n), .Y(n2899) );
 wddl_or U1901 ( .A(n2842), .A_n(n2842_n), .B(n2901), .B_n(n2901_n), .Y_n(n2880_n), .Y(n2880) );
 wddl_or U1902 ( .A(n2902), .A_n(n2902_n), .B(n2903), .B_n(n2903_n), .Y_n(n2901_n), .Y(n2901) );
 wddl_and U1903 ( .A(n2594), .A_n(n2594_n), .B(n2641), .B_n(n2641_n), .Y_n(n2903_n), .Y(n2903) );
 wddl_and U1904 ( .A(n2649), .A_n(n2649_n), .B(n2904), .B_n(n2904_n), .Y_n(n2902_n), .Y(n2902) );
 wddl_or U1905 ( .A(n2731), .A_n(n2731_n), .B(n2807), .B_n(n2807_n), .Y_n(n2878_n), .Y(n2878) );
 wddl_or U1906 ( .A(n2925), .A_n(n2925_n), .B(n2926), .B_n(n2926_n), .Y_n(n2807_n), .Y(n2807) );
 wddl_or U1907 ( .A(n2927), .A_n(n2927_n), .B(n2928), .B_n(n2928_n), .Y_n(n2926_n), .Y(n2926) );
 wddl_or U1908 ( .A(n2929), .A_n(n2929_n), .B(n2930), .B_n(n2930_n), .Y_n(n2928_n), .Y(n2928) );
 wddl_and U1909 ( .A(n2552), .A_n(n2552_n), .B(n2895), .B_n(n2895_n), .Y_n(n2930_n), .Y(n2930) );
 wddl_and U1910 ( .A(n2770), .A_n(n2770_n), .B(n2670), .B_n(n2670_n), .Y_n(n2929_n), .Y(n2929) );
 wddl_or U1911 ( .A(n2931), .A_n(n2931_n), .B(n2932), .B_n(n2932_n), .Y_n(n2927_n), .Y(n2927) );
 wddl_or U1912 ( .A(n2933), .A_n(n2933_n), .B(n2934), .B_n(n2934_n), .Y_n(n2932_n), .Y(n2932) );
 wddl_and U1913 ( .A(n2648), .A_n(n2648_n), .B(n2565), .B_n(n2565_n), .Y_n(n2934_n), .Y(n2934) );
 wddl_and U1914 ( .A(n2680), .A_n(n2680_n), .B(n2654), .B_n(n2654_n), .Y_n(n2931_n), .Y(n2931) );
 wddl_or U1915 ( .A(n2935), .A_n(n2935_n), .B(n2936), .B_n(n2936_n), .Y_n(n2925_n), .Y(n2925) );
 wddl_or U1916 ( .A(n2937), .A_n(n2937_n), .B(n2938), .B_n(n2938_n), .Y_n(n2936_n), .Y(n2936) );
 wddl_and U1917 ( .A(n2616), .A_n(n2616_n), .B(n2578), .B_n(n2578_n), .Y_n(n2938_n), .Y(n2938) );
 wddl_and U1918 ( .A(n2583), .A_n(n2583_n), .B(n2939), .B_n(n2939_n), .Y_n(n2937_n), .Y(n2937) );
 wddl_or U1919 ( .A(n2940), .A_n(n2940_n), .B(n2941), .B_n(n2941_n), .Y_n(n2935_n), .Y(n2935) );
 wddl_or U1920 ( .A(n2942), .A_n(n2942_n), .B(n2943), .B_n(n2943_n), .Y_n(n2941_n), .Y(n2941) );
 wddl_and U1921 ( .A(n2605), .A_n(n2605_n), .B(n2944), .B_n(n2944_n), .Y_n(n2943_n), .Y(n2943) );
 wddl_or U1922 ( .A(n2796), .A_n(n2796_n), .B(n2664), .B_n(n2664_n), .Y_n(n2944_n), .Y(n2944) );
 wddl_and U1923 ( .A(n2609), .A_n(n2609_n), .B(n2945), .B_n(n2945_n), .Y_n(n2942_n), .Y(n2942) );
 wddl_or U1924 ( .A(n2590), .A_n(n2590_n), .B(n2904), .B_n(n2904_n), .Y_n(n2945_n), .Y(n2945) );
 wddl_and U1925 ( .A(n2599), .A_n(n2599_n), .B(n2946), .B_n(n2946_n), .Y_n(n2940_n), .Y(n2940) );
 wddl_or U1926 ( .A(n2644), .A_n(n2644_n), .B(n2862), .B_n(n2862_n), .Y_n(n2946_n), .Y(n2946) );
 wddl_or U1927 ( .A(n2727), .A_n(n2727_n), .B(n2728), .B_n(n2728_n), .Y_n(d_n[7]), .Y(d[7]) );
 wddl_or U1928 ( .A(n2729), .A_n(n2729_n), .B(n2730), .B_n(n2730_n), .Y_n(n2728_n), .Y(n2728) );
 wddl_or U1929 ( .A(n2731), .A_n(n2731_n), .B(n2732), .B_n(n2732_n), .Y_n(n2730_n), .Y(n2730) );
 wddl_or U1930 ( .A(n2733), .A_n(n2733_n), .B(n2734), .B_n(n2734_n), .Y_n(n2732_n), .Y(n2732) );
 wddl_or U1931 ( .A(n2735), .A_n(n2735_n), .B(n2736), .B_n(n2736_n), .Y_n(n2733_n), .Y(n2733) );
 wddl_or U1932 ( .A(n2737), .A_n(n2737_n), .B(n2738), .B_n(n2738_n), .Y_n(n2736_n), .Y(n2736) );
 wddl_or U1933 ( .A(n2739), .A_n(n2739_n), .B(n2740), .B_n(n2740_n), .Y_n(n2738_n), .Y(n2738) );
 wddl_and U1934 ( .A(n2643), .A_n(n2643_n), .B(n2742), .B_n(n2742_n), .Y_n(n2740_n), .Y(n2740) );
 wddl_or U1935 ( .A(n2596), .A_n(n2596_n), .B(n2696), .B_n(n2696_n), .Y_n(n2742_n), .Y(n2742) );
 wddl_and U1936 ( .A(n2744), .A_n(n2744_n), .B(n2745), .B_n(n2745_n), .Y_n(n2739_n), .Y(n2739) );
 wddl_and U1937 ( .A(n2746), .A_n(n2746_n), .B(n2747), .B_n(n2747_n), .Y_n(n2737_n), .Y(n2737) );
 wddl_or U1938 ( .A(n2616), .A_n(n2616_n), .B(n2749), .B_n(n2749_n), .Y_n(n2747_n), .Y(n2747) );
 wddl_or U1939 ( .A(n2750), .A_n(n2750_n), .B(n2751), .B_n(n2751_n), .Y_n(n2735_n), .Y(n2735) );
 wddl_or U1940 ( .A(n2752), .A_n(n2752_n), .B(n2753), .B_n(n2753_n), .Y_n(n2751_n), .Y(n2751) );
 wddl_or U1941 ( .A(n2754), .A_n(n2754_n), .B(n2755), .B_n(n2755_n), .Y_n(n2753_n), .Y(n2753) );
 wddl_and U1942 ( .A(n2684), .A_n(n2684_n), .B(n2583), .B_n(n2583_n), .Y_n(n2755_n), .Y(n2755) );
 wddl_and U1943 ( .A(n2533), .A_n(n2533_n), .B(n2759), .B_n(n2759_n), .Y_n(n2754_n), .Y(n2754) );
 wddl_and U1944 ( .A(n2649), .A_n(n2649_n), .B(n2761), .B_n(n2761_n), .Y_n(n2752_n), .Y(n2752) );
 wddl_and U1945 ( .A(n2575), .A_n(n2575_n), .B(n2763), .B_n(n2763_n), .Y_n(n2750_n), .Y(n2750) );
 wddl_or U1946 ( .A(n2636), .A_n(n2636_n), .B(n2765), .B_n(n2765_n), .Y_n(n2763_n), .Y(n2763) );
 wddl_or U1947 ( .A(n2947), .A_n(n2947_n), .B(n2948), .B_n(n2948_n), .Y_n(n2731_n), .Y(n2731) );
 wddl_or U1948 ( .A(n2949), .A_n(n2949_n), .B(n2950), .B_n(n2950_n), .Y_n(n2948_n), .Y(n2948) );
 wddl_or U1949 ( .A(n2951), .A_n(n2951_n), .B(n2952), .B_n(n2952_n), .Y_n(n2950_n), .Y(n2950) );
 wddl_and U1950 ( .A(n2544), .A_n(n2544_n), .B(n2618), .B_n(n2618_n), .Y_n(n2952_n), .Y(n2952) );
 wddl_or U1951 ( .A(n2953), .A_n(n2953_n), .B(n2954), .B_n(n2954_n), .Y_n(n2949_n), .Y(n2949) );
 wddl_or U1952 ( .A(n2955), .A_n(n2955_n), .B(n2956), .B_n(n2956_n), .Y_n(n2954_n), .Y(n2954) );
 wddl_and U1953 ( .A(n2555), .A_n(n2555_n), .B(n2698), .B_n(n2698_n), .Y_n(n2956_n), .Y(n2956) );
 wddl_and U1954 ( .A(n2645), .A_n(n2645_n), .B(n2653), .B_n(n2653_n), .Y_n(n2955_n), .Y(n2955) );
 wddl_and U1955 ( .A(n2625), .A_n(n2625_n), .B(n2574), .B_n(n2574_n), .Y_n(n2953_n), .Y(n2953) );
 wddl_or U1956 ( .A(n2957), .A_n(n2957_n), .B(n2958), .B_n(n2958_n), .Y_n(n2947_n), .Y(n2947) );
 wddl_or U1957 ( .A(n2959), .A_n(n2959_n), .B(n2960), .B_n(n2960_n), .Y_n(n2958_n), .Y(n2958) );
 wddl_or U1958 ( .A(n2961), .A_n(n2961_n), .B(n2962), .B_n(n2962_n), .Y_n(n2960_n), .Y(n2960) );
 wddl_and U1959 ( .A(n2663), .A_n(n2663_n), .B(n2875), .B_n(n2875_n), .Y_n(n2962_n), .Y(n2962) );
 wddl_and U1960 ( .A(n2694), .A_n(n2694_n), .B(n2691), .B_n(n2691_n), .Y_n(n2961_n), .Y(n2961) );
 wddl_and U1961 ( .A(n2589), .A_n(n2589_n), .B(n2841), .B_n(n2841_n), .Y_n(n2959_n), .Y(n2959) );
 wddl_or U1962 ( .A(n2963), .A_n(n2963_n), .B(n2964), .B_n(n2964_n), .Y_n(n2957_n), .Y(n2957) );
 wddl_or U1963 ( .A(n2965), .A_n(n2965_n), .B(n2966), .B_n(n2966_n), .Y_n(n2964_n), .Y(n2964) );
 wddl_and U1964 ( .A(n2638), .A_n(n2638_n), .B(n2967), .B_n(n2967_n), .Y_n(n2966_n), .Y(n2966) );
 wddl_and U1965 ( .A(n2707), .A_n(n2707_n), .B(n2968), .B_n(n2968_n), .Y_n(n2965_n), .Y(n2965) );
 wddl_or U1966 ( .A(n2675), .A_n(n2675_n), .B(n2608), .B_n(n2608_n), .Y_n(n2968_n), .Y(n2968) );
 wddl_and U1967 ( .A(n2603), .A_n(n2603_n), .B(n2969), .B_n(n2969_n), .Y_n(n2963_n), .Y(n2963) );
 wddl_or U1968 ( .A(n2766), .A_n(n2766_n), .B(n2767), .B_n(n2767_n), .Y_n(n2729_n), .Y(n2729) );
 wddl_or U1969 ( .A(n2768), .A_n(n2768_n), .B(n2769), .B_n(n2769_n), .Y_n(n2767_n), .Y(n2767) );
 wddl_and U1970 ( .A(n2624), .A_n(n2624_n), .B(n2604), .B_n(n2604_n), .Y_n(n2769_n), .Y(n2769) );
 wddl_and U1971 ( .A(n2674), .A_n(n2674_n), .B(n2630), .B_n(n2630_n), .Y_n(n2768_n), .Y(n2768) );
 wddl_or U1972 ( .A(n2812), .A_n(n2812_n), .B(n2813), .B_n(n2813_n), .Y_n(n2727_n), .Y(n2727) );
 wddl_or U1973 ( .A(n2814), .A_n(n2814_n), .B(n2815), .B_n(n2815_n), .Y_n(n2813_n), .Y(n2813) );
 wddl_or U1974 ( .A(n2816), .A_n(n2816_n), .B(n2817), .B_n(n2817_n), .Y_n(n2815_n), .Y(n2815) );
 wddl_or U1975 ( .A(n2818), .A_n(n2818_n), .B(n2819), .B_n(n2819_n), .Y_n(n2817_n), .Y(n2817) );
 wddl_or U1976 ( .A(n2820), .A_n(n2820_n), .B(n2821), .B_n(n2821_n), .Y_n(n2819_n), .Y(n2819) );
 wddl_and U1977 ( .A(n2600), .A_n(n2600_n), .B(n2639), .B_n(n2639_n), .Y_n(n2820_n), .Y(n2820) );
 wddl_and U1978 ( .A(n2759), .A_n(n2759_n), .B(n2594), .B_n(n2594_n), .Y_n(n2818_n), .Y(n2818) );
 wddl_or U1979 ( .A(n2823), .A_n(n2823_n), .B(n2824), .B_n(n2824_n), .Y_n(n2814_n), .Y(n2814) );
 wddl_or U1980 ( .A(n2825), .A_n(n2825_n), .B(n2826), .B_n(n2826_n), .Y_n(n2824_n), .Y(n2824) );
 wddl_or U1981 ( .A(n2827), .A_n(n2827_n), .B(n2828), .B_n(n2828_n), .Y_n(n2826_n), .Y(n2826) );
 wddl_and U1982 ( .A(n2591), .A_n(n2591_n), .B(n2700), .B_n(n2700_n), .Y_n(n2828_n), .Y(n2828) );
 wddl_and U1983 ( .A(n2829), .A_n(n2829_n), .B(n2540), .B_n(n2540_n), .Y_n(n2827_n), .Y(n2827) );
 wddl_and U1984 ( .A(n2626), .A_n(n2626_n), .B(n2558), .B_n(n2558_n), .Y_n(n2825_n), .Y(n2825) );
 wddl_or U1985 ( .A(n2831), .A_n(n2831_n), .B(n2832), .B_n(n2832_n), .Y_n(n2823_n), .Y(n2823) );
 wddl_or U1986 ( .A(n2833), .A_n(n2833_n), .B(n2834), .B_n(n2834_n), .Y_n(n2832_n), .Y(n2832) );
 wddl_and U1987 ( .A(n2835), .A_n(n2835_n), .B(n2666), .B_n(n2666_n), .Y_n(n2834_n), .Y(n2834) );
 wddl_and U1988 ( .A(n2630), .A_n(n2630_n), .B(n2836), .B_n(n2836_n), .Y_n(n2833_n), .Y(n2833) );
 wddl_or U1989 ( .A(n2837), .A_n(n2837_n), .B(n2838), .B_n(n2838_n), .Y_n(n2831_n), .Y(n2831) );
 wddl_and U1990 ( .A(n2800), .A_n(n2800_n), .B(n2839), .B_n(n2839_n), .Y_n(n2838_n), .Y(n2838) );
 wddl_and U1991 ( .A(n2668), .A_n(n2668_n), .B(n2840), .B_n(n2840_n), .Y_n(n2837_n), .Y(n2837) );
 wddl_or U1992 ( .A(n2601), .A_n(n2601_n), .B(n2841), .B_n(n2841_n), .Y_n(n2840_n), .Y(n2840) );
 wddl_or U1993 ( .A(n2673), .A_n(n2673_n), .B(n2633), .B_n(n2633_n), .Y_n(n2841_n), .Y(n2841) );
 wddl_or U1994 ( .A(n2842), .A_n(n2842_n), .B(n2843), .B_n(n2843_n), .Y_n(n2812_n), .Y(n2812) );
 wddl_or U1995 ( .A(n2905), .A_n(n2905_n), .B(n2906), .B_n(n2906_n), .Y_n(n2842_n), .Y(n2842) );
 wddl_or U1996 ( .A(n2907), .A_n(n2907_n), .B(n2908), .B_n(n2908_n), .Y_n(n2906_n), .Y(n2906) );
 wddl_or U1997 ( .A(n2909), .A_n(n2909_n), .B(n2910), .B_n(n2910_n), .Y_n(n2908_n), .Y(n2908) );
 wddl_and U1998 ( .A(n2578), .A_n(n2578_n), .B(n2911), .B_n(n2911_n), .Y_n(n2910_n), .Y(n2910) );
 wddl_and U1999 ( .A(n2595), .A_n(n2595_n), .B(n2559), .B_n(n2559_n), .Y_n(n2909_n), .Y(n2909) );
 wddl_and U2000 ( .A(n2634), .A_n(n2634_n), .B(n2912), .B_n(n2912_n), .Y_n(n2907_n), .Y(n2907) );
 wddl_or U2001 ( .A(n2561), .A_n(n2561_n), .B(n2679), .B_n(n2679_n), .Y_n(n2912_n), .Y(n2912) );
 wddl_or U2002 ( .A(n2913), .A_n(n2913_n), .B(n2914), .B_n(n2914_n), .Y_n(n2905_n), .Y(n2905) );
 wddl_or U2003 ( .A(n2915), .A_n(n2915_n), .B(n2916), .B_n(n2916_n), .Y_n(n2914_n), .Y(n2914) );
 wddl_and U2004 ( .A(n2599), .A_n(n2599_n), .B(n2917), .B_n(n2917_n), .Y_n(n2916_n), .Y(n2916) );
 wddl_or U2005 ( .A(n2590), .A_n(n2590_n), .B(n2918), .B_n(n2918_n), .Y_n(n2917_n), .Y(n2917) );
 wddl_or U2006 ( .A(n2566), .A_n(n2566_n), .B(n2606), .B_n(n2606_n), .Y_n(n2918_n), .Y(n2918) );
 wddl_and U2007 ( .A(n2623), .A_n(n2623_n), .B(n2919), .B_n(n2919_n), .Y_n(n2915_n), .Y(n2915) );
 wddl_or U2008 ( .A(n2705), .A_n(n2705_n), .B(n2920), .B_n(n2920_n), .Y_n(n2919_n), .Y(n2919) );
 wddl_or U2009 ( .A(n2579), .A_n(n2579_n), .B(n2643), .B_n(n2643_n), .Y_n(n2920_n), .Y(n2920) );
 wddl_or U2010 ( .A(n2921), .A_n(n2921_n), .B(n2922), .B_n(n2922_n), .Y_n(n2913_n), .Y(n2913) );
 wddl_and U2011 ( .A(n2650), .A_n(n2650_n), .B(n2923), .B_n(n2923_n), .Y_n(n2922_n), .Y(n2922) );
 wddl_or U2012 ( .A(n2631), .A_n(n2631_n), .B(n2708), .B_n(n2708_n), .Y_n(n2923_n), .Y(n2923) );
 wddl_and U2013 ( .A(n2684), .A_n(n2684_n), .B(n2924), .B_n(n2924_n), .Y_n(n2921_n), .Y(n2921) );
 wddl_or U2014 ( .A(n2748), .A_n(n2748_n), .B(n2674), .B_n(n2674_n), .Y_n(n2924_n), .Y(n2924) );
 wddl_or U2015 ( .A(n2844), .A_n(n2844_n), .B(n2970), .B_n(n2970_n), .Y_n(d_n[3]), .Y(d[3]) );
 wddl_or U2016 ( .A(n2971), .A_n(n2971_n), .B(n2972), .B_n(n2972_n), .Y_n(n2970_n), .Y(n2970) );
 wddl_or U2017 ( .A(n2973), .A_n(n2973_n), .B(n2974), .B_n(n2974_n), .Y_n(n2972_n), .Y(n2972) );
 wddl_or U2018 ( .A(n2975), .A_n(n2975_n), .B(n2976), .B_n(n2976_n), .Y_n(n2974_n), .Y(n2974) );
 wddl_or U2019 ( .A(n2977), .A_n(n2977_n), .B(n2978), .B_n(n2978_n), .Y_n(n2976_n), .Y(n2976) );
 wddl_and U2020 ( .A(n2874), .A_n(n2874_n), .B(n2979), .B_n(n2979_n), .Y_n(n2978_n), .Y(n2978) );
 wddl_and U2021 ( .A(n2699), .A_n(n2699_n), .B(n2576), .B_n(n2576_n), .Y_n(n2977_n), .Y(n2977) );
 wddl_and U2022 ( .A(n2709), .A_n(n2709_n), .B(n2651), .B_n(n2651_n), .Y_n(n2975_n), .Y(n2975) );
 wddl_or U2023 ( .A(n2980), .A_n(n2980_n), .B(n2981), .B_n(n2981_n), .Y_n(n2971_n), .Y(n2971) );
 wddl_or U2024 ( .A(n2982), .A_n(n2982_n), .B(n2983), .B_n(n2983_n), .Y_n(n2981_n), .Y(n2981) );
 wddl_or U2025 ( .A(n3330), .A_n(n3330_n), .B(n3331), .B_n(n3331_n), .Y_n(n2983_n), .Y(n2983) );
 wddl_or U2026 ( .A(n3332), .A_n(n3332_n), .B(n3333), .B_n(n3333_n), .Y_n(n3331_n), .Y(n3331) );
 wddl_or U2027 ( .A(n3334), .A_n(n3334_n), .B(n3335), .B_n(n3335_n), .Y_n(n3333_n), .Y(n3333) );
 wddl_or U2028 ( .A(n3224), .A_n(n3224_n), .B(n2821), .B_n(n2821_n), .Y_n(n3335_n), .Y(n3335) );
 wddl_and U2029 ( .A(n2686), .A_n(n2686_n), .B(n2620), .B_n(n2620_n), .Y_n(n2821_n), .Y(n2821) );
 wddl_and U2030 ( .A(n2581), .A_n(n2581_n), .B(n2869), .B_n(n2869_n), .Y_n(n3334_n), .Y(n3334) );
 wddl_or U2031 ( .A(n2772), .A_n(n2772_n), .B(n2621), .B_n(n2621_n), .Y_n(n2869_n), .Y(n2869) );
 wddl_and U2032 ( .A(n2601), .A_n(n2601_n), .B(n2888), .B_n(n2888_n), .Y_n(n3332_n), .Y(n3332) );
 wddl_or U2033 ( .A(n3336), .A_n(n3336_n), .B(n3337), .B_n(n3337_n), .Y_n(n3330_n), .Y(n3330) );
 wddl_or U2034 ( .A(n3338), .A_n(n3338_n), .B(n3339), .B_n(n3339_n), .Y_n(n3337_n), .Y(n3337) );
 wddl_and U2035 ( .A(n2606), .A_n(n2606_n), .B(n2520), .B_n(n2520_n), .Y_n(n3339_n), .Y(n3339) );
 wddl_and U2036 ( .A(n2695), .A_n(n2695_n), .B(n3072), .B_n(n3072_n), .Y_n(n3338_n), .Y(n3338) );
 wddl_or U2037 ( .A(n3340), .A_n(n3340_n), .B(n3341), .B_n(n3341_n), .Y_n(n3336_n), .Y(n3336) );
 wddl_and U2038 ( .A(n2705), .A_n(n2705_n), .B(n3342), .B_n(n3342_n), .Y_n(n3341_n), .Y(n3341) );
 wddl_or U2039 ( .A(n2623), .A_n(n2623_n), .B(n2619), .B_n(n2619_n), .Y_n(n3342_n), .Y(n3342) );
 wddl_and U2040 ( .A(n2661), .A_n(n2661_n), .B(n3343), .B_n(n3343_n), .Y_n(n3340_n), .Y(n3340) );
 wddl_or U2041 ( .A(n2530), .A_n(n2530_n), .B(n2904), .B_n(n2904_n), .Y_n(n3343_n), .Y(n3343) );
 wddl_or U2042 ( .A(n2984), .A_n(n2984_n), .B(n2985), .B_n(n2985_n), .Y_n(n2982_n), .Y(n2982) );
 wddl_or U2043 ( .A(n2986), .A_n(n2986_n), .B(n2987), .B_n(n2987_n), .Y_n(n2985_n), .Y(n2985) );
 wddl_and U2044 ( .A(n2623), .A_n(n2623_n), .B(n2988), .B_n(n2988_n), .Y_n(n2987_n), .Y(n2987) );
 wddl_or U2045 ( .A(n2628), .A_n(n2628_n), .B(n2558), .B_n(n2558_n), .Y_n(n2988_n), .Y(n2988) );
 wddl_and U2046 ( .A(n2565), .A_n(n2565_n), .B(n2989), .B_n(n2989_n), .Y_n(n2986_n), .Y(n2986) );
 wddl_or U2047 ( .A(n2615), .A_n(n2615_n), .B(n2990), .B_n(n2990_n), .Y_n(n2989_n), .Y(n2989) );
 wddl_or U2048 ( .A(n2991), .A_n(n2991_n), .B(n2992), .B_n(n2992_n), .Y_n(n2984_n), .Y(n2984) );
 wddl_or U2049 ( .A(n2993), .A_n(n2993_n), .B(n2994), .B_n(n2994_n), .Y_n(n2992_n), .Y(n2992) );
 wddl_and U2050 ( .A(n2522), .A_n(n2522_n), .B(n2656), .B_n(n2656_n), .Y_n(n2994_n), .Y(n2994) );
 wddl_and U2051 ( .A(n2689), .A_n(n2689_n), .B(n2996), .B_n(n2996_n), .Y_n(n2993_n), .Y(n2993) );
 wddl_or U2052 ( .A(n2600), .A_n(n2600_n), .B(n2693), .B_n(n2693_n), .Y_n(n2996_n), .Y(n2996) );
 wddl_or U2053 ( .A(n2997), .A_n(n2997_n), .B(n2998), .B_n(n2998_n), .Y_n(n2991_n), .Y(n2991) );
 wddl_or U2054 ( .A(n2999), .A_n(n2999_n), .B(n3000), .B_n(n3000_n), .Y_n(n2998_n), .Y(n2998) );
 wddl_and U2055 ( .A(n2741), .A_n(n2741_n), .B(n2571), .B_n(n2571_n), .Y_n(n3000_n), .Y(n3000) );
 wddl_and U2056 ( .A(n2585), .A_n(n2585_n), .B(n2640), .B_n(n2640_n), .Y_n(n2999_n), .Y(n2999) );
 wddl_and U2057 ( .A(n2590), .A_n(n2590_n), .B(n2550), .B_n(n2550_n), .Y_n(n2997_n), .Y(n2997) );
 wddl_or U2058 ( .A(n3001), .A_n(n3001_n), .B(n3002), .B_n(n3002_n), .Y_n(n2844_n), .Y(n2844) );
 wddl_or U2059 ( .A(n3003), .A_n(n3003_n), .B(n3004), .B_n(n3004_n), .Y_n(n3002_n), .Y(n3002) );
 wddl_or U2060 ( .A(n3308), .A_n(n3308_n), .B(n3309), .B_n(n3309_n), .Y_n(n3004_n), .Y(n3004) );
 wddl_or U2061 ( .A(n3310), .A_n(n3310_n), .B(n3311), .B_n(n3311_n), .Y_n(n3309_n), .Y(n3309) );
 wddl_or U2062 ( .A(n3312), .A_n(n3312_n), .B(n3313), .B_n(n3313_n), .Y_n(n3311_n), .Y(n3311) );
 wddl_or U2063 ( .A(n3314), .A_n(n3314_n), .B(n3315), .B_n(n3315_n), .Y_n(n3313_n), .Y(n3313) );
 wddl_and U2064 ( .A(n2552), .A_n(n2552_n), .B(n2598), .B_n(n2598_n), .Y_n(n3315_n), .Y(n3315) );
 wddl_and U2065 ( .A(n2700), .A_n(n2700_n), .B(n2797), .B_n(n2797_n), .Y_n(n3314_n), .Y(n3314) );
 wddl_and U2066 ( .A(n2676), .A_n(n2676_n), .B(n2680), .B_n(n2680_n), .Y_n(n3312_n), .Y(n3312) );
 wddl_or U2067 ( .A(n3316), .A_n(n3316_n), .B(n3317), .B_n(n3317_n), .Y_n(n3310_n), .Y(n3310) );
 wddl_or U2068 ( .A(n3318), .A_n(n3318_n), .B(n3319), .B_n(n3319_n), .Y_n(n3317_n), .Y(n3317) );
 wddl_and U2069 ( .A(n2608), .A_n(n2608_n), .B(n2671), .B_n(n2671_n), .Y_n(n3319_n), .Y(n3319) );
 wddl_and U2070 ( .A(n2705), .A_n(n2705_n), .B(n2538), .B_n(n2538_n), .Y_n(n3318_n), .Y(n3318) );
 wddl_and U2071 ( .A(n2770), .A_n(n2770_n), .B(n2566), .B_n(n2566_n), .Y_n(n3316_n), .Y(n3316) );
 wddl_or U2072 ( .A(n3320), .A_n(n3320_n), .B(n3321), .B_n(n3321_n), .Y_n(n3308_n), .Y(n3308) );
 wddl_or U2073 ( .A(n3322), .A_n(n3322_n), .B(n3323), .B_n(n3323_n), .Y_n(n3321_n), .Y(n3321) );
 wddl_or U2074 ( .A(n3324), .A_n(n3324_n), .B(n3325), .B_n(n3325_n), .Y_n(n3323_n), .Y(n3323) );
 wddl_and U2075 ( .A(n2650), .A_n(n2650_n), .B(n2581), .B_n(n2581_n), .Y_n(n3325_n), .Y(n3325) );
 wddl_and U2076 ( .A(n2656), .A_n(n2656_n), .B(n2904), .B_n(n2904_n), .Y_n(n3324_n), .Y(n3324) );
 wddl_or U2077 ( .A(n2703), .A_n(n2703_n), .B(n2670), .B_n(n2670_n), .Y_n(n2904_n), .Y(n2904) );
 wddl_and U2078 ( .A(n2630), .A_n(n2630_n), .B(n2765), .B_n(n2765_n), .Y_n(n3322_n), .Y(n3322) );
 wddl_or U2079 ( .A(n3326), .A_n(n3326_n), .B(n3327), .B_n(n3327_n), .Y_n(n3320_n), .Y(n3320) );
 wddl_or U2080 ( .A(n3183), .A_n(n3183_n), .B(n3328), .B_n(n3328_n), .Y_n(n3327_n), .Y(n3327) );
 wddl_and U2081 ( .A(n2830), .A_n(n2830_n), .B(n2990), .B_n(n2990_n), .Y_n(n3328_n), .Y(n3328) );
 wddl_and U2082 ( .A(n2594), .A_n(n2594_n), .B(n3329), .B_n(n3329_n), .Y_n(n3326_n), .Y(n3326) );
 wddl_or U2083 ( .A(n2581), .A_n(n2581_n), .B(n2641), .B_n(n2641_n), .Y_n(n3329_n), .Y(n3329) );
 wddl_or U2084 ( .A(n3005), .A_n(n3005_n), .B(n3006), .B_n(n3006_n), .Y_n(n3003_n), .Y(n3003) );
 wddl_or U2085 ( .A(n3007), .A_n(n3007_n), .B(n3008), .B_n(n3008_n), .Y_n(n3006_n), .Y(n3006) );
 wddl_or U2086 ( .A(n3009), .A_n(n3009_n), .B(n3010), .B_n(n3010_n), .Y_n(n3008_n), .Y(n3008) );
 wddl_or U2087 ( .A(n3011), .A_n(n3011_n), .B(n3012), .B_n(n3012_n), .Y_n(n3010_n), .Y(n3010) );
 wddl_and U2088 ( .A(n2631), .A_n(n2631_n), .B(n2694), .B_n(n2694_n), .Y_n(n3012_n), .Y(n3012) );
 wddl_and U2089 ( .A(n2578), .A_n(n2578_n), .B(n3013), .B_n(n3013_n), .Y_n(n3011_n), .Y(n3011) );
 wddl_or U2090 ( .A(n2660), .A_n(n2660_n), .B(n3014), .B_n(n3014_n), .Y_n(n3013_n), .Y(n3013) );
 wddl_or U2091 ( .A(n2758), .A_n(n2758_n), .B(n2663), .B_n(n2663_n), .Y_n(n3014_n), .Y(n3014) );
 wddl_and U2092 ( .A(n2644), .A_n(n2644_n), .B(n3015), .B_n(n3015_n), .Y_n(n3009_n), .Y(n3009) );
 wddl_or U2093 ( .A(n3016), .A_n(n3016_n), .B(n3017), .B_n(n3017_n), .Y_n(n3007_n), .Y(n3007) );
 wddl_or U2094 ( .A(n3018), .A_n(n3018_n), .B(n3019), .B_n(n3019_n), .Y_n(n3017_n), .Y(n3017) );
 wddl_and U2095 ( .A(n2611), .A_n(n2611_n), .B(n3020), .B_n(n3020_n), .Y_n(n3019_n), .Y(n3019) );
 wddl_or U2096 ( .A(n2685), .A_n(n2685_n), .B(n2646), .B_n(n2646_n), .Y_n(n3020_n), .Y(n3020) );
 wddl_and U2097 ( .A(n2573), .A_n(n2573_n), .B(n3021), .B_n(n3021_n), .Y_n(n3018_n), .Y(n3018) );
 wddl_or U2098 ( .A(n2546), .A_n(n2546_n), .B(n2648), .B_n(n2648_n), .Y_n(n3021_n), .Y(n3021) );
 wddl_and U2099 ( .A(n2569), .A_n(n2569_n), .B(n3022), .B_n(n3022_n), .Y_n(n3016_n), .Y(n3016) );
 wddl_or U2100 ( .A(n2804), .A_n(n2804_n), .B(n2689), .B_n(n2689_n), .Y_n(n3022_n), .Y(n3022) );
 wddl_or U2101 ( .A(n3023), .A_n(n3023_n), .B(n3024), .B_n(n3024_n), .Y_n(n3001_n), .Y(n3001) );
 wddl_or U2102 ( .A(n3025), .A_n(n3025_n), .B(n3026), .B_n(n3026_n), .Y_n(n3024_n), .Y(n3024) );
 wddl_or U2103 ( .A(n2951), .A_n(n2951_n), .B(n3027), .B_n(n3027_n), .Y_n(n3026_n), .Y(n3026) );
 wddl_and U2104 ( .A(n2605), .A_n(n2605_n), .B(n2654), .B_n(n2654_n), .Y_n(n3027_n), .Y(n3027) );
 wddl_and U2105 ( .A(n2683), .A_n(n2683_n), .B(n2661), .B_n(n2661_n), .Y_n(n2951_n), .Y(n2951) );
 wddl_and U2106 ( .A(n2624), .A_n(n2624_n), .B(n2679), .B_n(n2679_n), .Y_n(n3025_n), .Y(n3025) );
 wddl_or U2107 ( .A(n3028), .A_n(n3028_n), .B(n3029), .B_n(n3029_n), .Y_n(d_n[2]), .Y(d[2]) );
 wddl_or U2108 ( .A(n3030), .A_n(n3030_n), .B(n3031), .B_n(n3031_n), .Y_n(n3029_n), .Y(n3029) );
 wddl_or U2109 ( .A(n3005), .A_n(n3005_n), .B(n3032), .B_n(n3032_n), .Y_n(n3031_n), .Y(n3031) );
 wddl_or U2110 ( .A(n3033), .A_n(n3033_n), .B(n3034), .B_n(n3034_n), .Y_n(n3032_n), .Y(n3032) );
 wddl_or U2111 ( .A(n3035), .A_n(n3035_n), .B(n3036), .B_n(n3036_n), .Y_n(n3034_n), .Y(n3034) );
 wddl_or U2112 ( .A(n3037), .A_n(n3037_n), .B(n3038), .B_n(n3038_n), .Y_n(n3036_n), .Y(n3036) );
 wddl_and U2113 ( .A(n2811), .A_n(n2811_n), .B(n2900), .B_n(n2900_n), .Y_n(n3038_n), .Y(n3038) );
 wddl_and U2114 ( .A(n2995), .A_n(n2995_n), .B(n2610), .B_n(n2610_n), .Y_n(n3037_n), .Y(n3037) );
 wddl_or U2115 ( .A(n3039), .A_n(n3039_n), .B(n3040), .B_n(n3040_n), .Y_n(n3035_n), .Y(n3035) );
 wddl_or U2116 ( .A(n3041), .A_n(n3041_n), .B(n3042), .B_n(n3042_n), .Y_n(n3040_n), .Y(n3040) );
 wddl_and U2117 ( .A(n2644), .A_n(n2644_n), .B(n2635), .B_n(n2635_n), .Y_n(n3042_n), .Y(n3042) );
 wddl_and U2118 ( .A(n2669), .A_n(n2669_n), .B(n2663), .B_n(n2663_n), .Y_n(n3041_n), .Y(n3041) );
 wddl_and U2119 ( .A(n2540), .A_n(n2540_n), .B(n2654), .B_n(n2654_n), .Y_n(n3039_n), .Y(n3039) );
 wddl_or U2120 ( .A(n3043), .A_n(n3043_n), .B(n3044), .B_n(n3044_n), .Y_n(n3033_n), .Y(n3033) );
 wddl_or U2121 ( .A(n3045), .A_n(n3045_n), .B(n3046), .B_n(n3046_n), .Y_n(n3044_n), .Y(n3044) );
 wddl_and U2122 ( .A(n2558), .A_n(n2558_n), .B(n3047), .B_n(n3047_n), .Y_n(n3046_n), .Y(n3046) );
 wddl_or U2123 ( .A(n3048), .A_n(n3048_n), .B(n2520), .B_n(n2520_n), .Y_n(n3047_n), .Y(n3047) );
 wddl_and U2124 ( .A(n2574), .A_n(n2574_n), .B(n3050), .B_n(n3050_n), .Y_n(n3045_n), .Y(n3045) );
 wddl_or U2125 ( .A(n2533), .A_n(n2533_n), .B(n2596), .B_n(n2596_n), .Y_n(n3050_n), .Y(n3050) );
 wddl_or U2126 ( .A(n3051), .A_n(n3051_n), .B(n3052), .B_n(n3052_n), .Y_n(n3043_n), .Y(n3043) );
 wddl_and U2127 ( .A(n2683), .A_n(n2683_n), .B(n2699), .B_n(n2699_n), .Y_n(n3052_n), .Y(n3052) );
 wddl_or U2128 ( .A(n3053), .A_n(n3053_n), .B(n3054), .B_n(n3054_n), .Y_n(n3005_n), .Y(n3005) );
 wddl_or U2129 ( .A(n3055), .A_n(n3055_n), .B(n3056), .B_n(n3056_n), .Y_n(n3054_n), .Y(n3054) );
 wddl_or U2130 ( .A(n3057), .A_n(n3057_n), .B(n3058), .B_n(n3058_n), .Y_n(n3056_n), .Y(n3056) );
 wddl_or U2131 ( .A(n3059), .A_n(n3059_n), .B(n3060), .B_n(n3060_n), .Y_n(n3058_n), .Y(n3058) );
 wddl_and U2132 ( .A(n2603), .A_n(n2603_n), .B(n2586), .B_n(n2586_n), .Y_n(n3060_n), .Y(n3060) );
 wddl_and U2133 ( .A(n2598), .A_n(n2598_n), .B(n2900), .B_n(n2900_n), .Y_n(n3057_n), .Y(n3057) );
 wddl_and U2134 ( .A(n2748), .A_n(n2748_n), .B(n2526), .B_n(n2526_n), .Y_n(n3055_n), .Y(n3055) );
 wddl_or U2135 ( .A(n3061), .A_n(n3061_n), .B(n3062), .B_n(n3062_n), .Y_n(n3053_n), .Y(n3053) );
 wddl_or U2136 ( .A(n3063), .A_n(n3063_n), .B(n3064), .B_n(n3064_n), .Y_n(n3062_n), .Y(n3062) );
 wddl_and U2137 ( .A(n2689), .A_n(n2689_n), .B(n3015), .B_n(n3015_n), .Y_n(n3064_n), .Y(n3064) );
 wddl_or U2138 ( .A(n2615), .A_n(n2615_n), .B(n2620), .B_n(n2620_n), .Y_n(n3015_n), .Y(n3015) );
 wddl_and U2139 ( .A(n2557), .A_n(n2557_n), .B(n3065), .B_n(n3065_n), .Y_n(n3063_n), .Y(n3063) );
 wddl_or U2140 ( .A(n3066), .A_n(n3066_n), .B(n3067), .B_n(n3067_n), .Y_n(n3061_n), .Y(n3061) );
 wddl_or U2141 ( .A(n3068), .A_n(n3068_n), .B(n3069), .B_n(n3069_n), .Y_n(n3067_n), .Y(n3067) );
 wddl_and U2142 ( .A(n2554), .A_n(n2554_n), .B(n3070), .B_n(n3070_n), .Y_n(n3069_n), .Y(n3069) );
 wddl_and U2143 ( .A(n2628), .A_n(n2628_n), .B(n3071), .B_n(n3071_n), .Y_n(n3068_n), .Y(n3068) );
 wddl_or U2144 ( .A(n2673), .A_n(n2673_n), .B(n2660), .B_n(n2660_n), .Y_n(n3071_n), .Y(n3071) );
 wddl_and U2145 ( .A(n2654), .A_n(n2654_n), .B(n3072), .B_n(n3072_n), .Y_n(n3066_n), .Y(n3066) );
 wddl_or U2146 ( .A(n2799), .A_n(n2799_n), .B(n2639), .B_n(n2639_n), .Y_n(n3072_n), .Y(n3072) );
 wddl_or U2147 ( .A(n2848), .A_n(n2848_n), .B(n2980), .B_n(n2980_n), .Y_n(n3030_n), .Y(n3030) );
 wddl_or U2148 ( .A(n3073), .A_n(n3073_n), .B(n3074), .B_n(n3074_n), .Y_n(n2980_n), .Y(n2980) );
 wddl_or U2149 ( .A(n3075), .A_n(n3075_n), .B(n3076), .B_n(n3076_n), .Y_n(n3074_n), .Y(n3074) );
 wddl_or U2150 ( .A(n3077), .A_n(n3077_n), .B(n3078), .B_n(n3078_n), .Y_n(n3076_n), .Y(n3076) );
 wddl_and U2151 ( .A(n2700), .A_n(n2700_n), .B(n2888), .B_n(n2888_n), .Y_n(n3078_n), .Y(n3078) );
 wddl_and U2152 ( .A(n2580), .A_n(n2580_n), .B(n2608), .B_n(n2608_n), .Y_n(n3077_n), .Y(n3077) );
 wddl_or U2153 ( .A(n2809), .A_n(n2809_n), .B(n3079), .B_n(n3079_n), .Y_n(n3075_n), .Y(n3075) );
 wddl_and U2154 ( .A(n2671), .A_n(n2671_n), .B(n3080), .B_n(n3080_n), .Y_n(n3079_n), .Y(n3079) );
 wddl_and U2155 ( .A(n2588), .A_n(n2588_n), .B(n2595), .B_n(n2595_n), .Y_n(n2809_n), .Y(n2809) );
 wddl_or U2156 ( .A(n3081), .A_n(n3081_n), .B(n3082), .B_n(n3082_n), .Y_n(n3073_n), .Y(n3073) );
 wddl_or U2157 ( .A(n3083), .A_n(n3083_n), .B(n3084), .B_n(n3084_n), .Y_n(n3082_n), .Y(n3082) );
 wddl_and U2158 ( .A(n2555), .A_n(n2555_n), .B(n3085), .B_n(n3085_n), .Y_n(n3084_n), .Y(n3084) );
 wddl_and U2159 ( .A(n2616), .A_n(n2616_n), .B(n3086), .B_n(n3086_n), .Y_n(n3083_n), .Y(n3083) );
 wddl_or U2160 ( .A(n2680), .A_n(n2680_n), .B(n2862), .B_n(n2862_n), .Y_n(n3086_n), .Y(n3086) );
 wddl_or U2161 ( .A(n3087), .A_n(n3087_n), .B(n3088), .B_n(n3088_n), .Y_n(n3081_n), .Y(n3081) );
 wddl_and U2162 ( .A(n2646), .A_n(n2646_n), .B(n3089), .B_n(n3089_n), .Y_n(n3088_n), .Y(n3088) );
 wddl_or U2163 ( .A(n2661), .A_n(n2661_n), .B(n2653), .B_n(n2653_n), .Y_n(n3089_n), .Y(n3089) );
 wddl_and U2164 ( .A(n2696), .A_n(n2696_n), .B(n3090), .B_n(n3090_n), .Y_n(n3087_n), .Y(n3087) );
 wddl_or U2165 ( .A(n2604), .A_n(n2604_n), .B(n2530), .B_n(n2530_n), .Y_n(n3090_n), .Y(n3090) );
 wddl_or U2166 ( .A(n3091), .A_n(n3091_n), .B(n3092), .B_n(n3092_n), .Y_n(n2848_n), .Y(n2848) );
 wddl_or U2167 ( .A(n3093), .A_n(n3093_n), .B(n3094), .B_n(n3094_n), .Y_n(n3092_n), .Y(n3092) );
 wddl_or U2168 ( .A(n3095), .A_n(n3095_n), .B(n3096), .B_n(n3096_n), .Y_n(n3094_n), .Y(n3094) );
 wddl_and U2169 ( .A(n2676), .A_n(n2676_n), .B(n2684), .B_n(n2684_n), .Y_n(n3096_n), .Y(n3096) );
 wddl_or U2170 ( .A(n3097), .A_n(n3097_n), .B(n3098), .B_n(n3098_n), .Y_n(n3093_n), .Y(n3093) );
 wddl_or U2171 ( .A(n2933), .A_n(n2933_n), .B(n3099), .B_n(n3099_n), .Y_n(n3098_n), .Y(n3098) );
 wddl_and U2172 ( .A(n2628), .A_n(n2628_n), .B(n2634), .B_n(n2634_n), .Y_n(n3099_n), .Y(n3099) );
 wddl_and U2173 ( .A(n2658), .A_n(n2658_n), .B(n2690), .B_n(n2690_n), .Y_n(n2933_n), .Y(n2933) );
 wddl_or U2174 ( .A(n3100), .A_n(n3100_n), .B(n3101), .B_n(n3101_n), .Y_n(n3091_n), .Y(n3091) );
 wddl_or U2175 ( .A(n3102), .A_n(n3102_n), .B(n3103), .B_n(n3103_n), .Y_n(n3101_n), .Y(n3101) );
 wddl_and U2176 ( .A(n2664), .A_n(n2664_n), .B(n3104), .B_n(n3104_n), .Y_n(n3103_n), .Y(n3103) );
 wddl_or U2177 ( .A(n2544), .A_n(n2544_n), .B(n2574), .B_n(n2574_n), .Y_n(n3104_n), .Y(n3104) );
 wddl_and U2178 ( .A(n2668), .A_n(n2668_n), .B(n3105), .B_n(n3105_n), .Y_n(n3102_n), .Y(n3102) );
 wddl_or U2179 ( .A(n2674), .A_n(n2674_n), .B(n2694), .B_n(n2694_n), .Y_n(n3105_n), .Y(n3105) );
 wddl_or U2180 ( .A(n3106), .A_n(n3106_n), .B(n3107), .B_n(n3107_n), .Y_n(n3100_n), .Y(n3100) );
 wddl_or U2181 ( .A(n3108), .A_n(n3108_n), .B(n3109), .B_n(n3109_n), .Y_n(n3107_n), .Y(n3107) );
 wddl_or U2182 ( .A(n3110), .A_n(n3110_n), .B(n3111), .B_n(n3111_n), .Y_n(n3109_n), .Y(n3109) );
 wddl_and U2183 ( .A(n2710), .A_n(n2710_n), .B(n3048), .B_n(n3048_n), .Y_n(n3111_n), .Y(n3111) );
 wddl_and U2184 ( .A(n2562), .A_n(n2562_n), .B(n2584), .B_n(n2584_n), .Y_n(n3110_n), .Y(n3110) );
 wddl_and U2185 ( .A(n2596), .A_n(n2596_n), .B(n3112), .B_n(n3112_n), .Y_n(n3108_n), .Y(n3108) );
 wddl_and U2186 ( .A(n2613), .A_n(n2613_n), .B(n3113), .B_n(n3113_n), .Y_n(n3106_n), .Y(n3106) );
 wddl_or U2187 ( .A(n2805), .A_n(n2805_n), .B(n2638), .B_n(n2638_n), .Y_n(n3113_n), .Y(n3113) );
 wddl_or U2188 ( .A(n3362), .A_n(n3362_n), .B(n3363), .B_n(n3363_n), .Y_n(n3028_n), .Y(n3028) );
 wddl_or U2189 ( .A(n2851), .A_n(n2851_n), .B(n3364), .B_n(n3364_n), .Y_n(n3363_n), .Y(n3363) );
 wddl_or U2190 ( .A(n2973), .A_n(n2973_n), .B(n3365), .B_n(n3365_n), .Y_n(n3364_n), .Y(n3364) );
 wddl_or U2191 ( .A(n3366), .A_n(n3366_n), .B(n3367), .B_n(n3367_n), .Y_n(n3365_n), .Y(n3365) );
 wddl_or U2192 ( .A(n3368), .A_n(n3368_n), .B(n3369), .B_n(n3369_n), .Y_n(n3367_n), .Y(n3367) );
 wddl_or U2193 ( .A(n3370), .A_n(n3370_n), .B(n3371), .B_n(n3371_n), .Y_n(n3369_n), .Y(n3369) );
 wddl_and U2194 ( .A(n2764), .A_n(n2764_n), .B(n2979), .B_n(n2979_n), .Y_n(n3371_n), .Y(n3371) );
 wddl_and U2195 ( .A(n2673), .A_n(n2673_n), .B(n2688), .B_n(n2688_n), .Y_n(n3370_n), .Y(n3370) );
 wddl_and U2196 ( .A(n2644), .A_n(n2644_n), .B(n2626), .B_n(n2626_n), .Y_n(n3368_n), .Y(n3368) );
 wddl_or U2197 ( .A(n3372), .A_n(n3372_n), .B(n3373), .B_n(n3373_n), .Y_n(n3366_n), .Y(n3366) );
 wddl_or U2198 ( .A(n3374), .A_n(n3374_n), .B(n3375), .B_n(n3375_n), .Y_n(n3373_n), .Y(n3373) );
 wddl_or U2199 ( .A(n3376), .A_n(n3376_n), .B(n3377), .B_n(n3377_n), .Y_n(n3375_n), .Y(n3375) );
 wddl_and U2200 ( .A(n2586), .A_n(n2586_n), .B(n3145), .B_n(n3145_n), .Y_n(n3377_n), .Y(n3377) );
 wddl_and U2201 ( .A(n2759), .A_n(n2759_n), .B(n3378), .B_n(n3378_n), .Y_n(n3376_n), .Y(n3376) );
 wddl_or U2202 ( .A(n2571), .A_n(n2571_n), .B(n2621), .B_n(n2621_n), .Y_n(n3378_n), .Y(n3378) );
 wddl_and U2203 ( .A(n2788), .A_n(n2788_n), .B(n3070), .B_n(n3070_n), .Y_n(n3374_n), .Y(n3374) );
 wddl_or U2204 ( .A(n2649), .A_n(n2649_n), .B(n2822), .B_n(n2822_n), .Y_n(n3070_n), .Y(n3070) );
 wddl_and U2205 ( .A(n2613), .A_n(n2613_n), .B(n3379), .B_n(n3379_n), .Y_n(n3372_n), .Y(n3372) );
 wddl_or U2206 ( .A(n2707), .A_n(n2707_n), .B(n2668), .B_n(n2668_n), .Y_n(n3379_n), .Y(n3379) );
 wddl_or U2207 ( .A(n3381), .A_n(n3381_n), .B(n3382), .B_n(n3382_n), .Y_n(n2973_n), .Y(n2973) );
 wddl_or U2208 ( .A(n3383), .A_n(n3383_n), .B(n3384), .B_n(n3384_n), .Y_n(n3382_n), .Y(n3382) );
 wddl_or U2209 ( .A(n3385), .A_n(n3385_n), .B(n3386), .B_n(n3386_n), .Y_n(n3384_n), .Y(n3384) );
 wddl_and U2210 ( .A(n2633), .A_n(n2633_n), .B(n3387), .B_n(n3387_n), .Y_n(n3386_n), .Y(n3386) );
 wddl_or U2211 ( .A(n2705), .A_n(n2705_n), .B(n2591), .B_n(n2591_n), .Y_n(n3387_n), .Y(n3387) );
 wddl_and U2212 ( .A(n2698), .A_n(n2698_n), .B(n3388), .B_n(n3388_n), .Y_n(n3385_n), .Y(n3385) );
 wddl_or U2213 ( .A(n2579), .A_n(n2579_n), .B(n2688), .B_n(n2688_n), .Y_n(n3388_n), .Y(n3388) );
 wddl_and U2214 ( .A(n2804), .A_n(n2804_n), .B(n3389), .B_n(n3389_n), .Y_n(n3383_n), .Y(n3383) );
 wddl_or U2215 ( .A(n2595), .A_n(n2595_n), .B(n2661), .B_n(n2661_n), .Y_n(n3389_n), .Y(n3389) );
 wddl_or U2216 ( .A(n3390), .A_n(n3390_n), .B(n3391), .B_n(n3391_n), .Y_n(n3381_n), .Y(n3381) );
 wddl_or U2217 ( .A(n3392), .A_n(n3392_n), .B(n3393), .B_n(n3393_n), .Y_n(n3391_n), .Y(n3391) );
 wddl_or U2218 ( .A(n3394), .A_n(n3394_n), .B(n3395), .B_n(n3395_n), .Y_n(n3393_n), .Y(n3393) );
 wddl_and U2219 ( .A(n2643), .A_n(n2643_n), .B(n2693), .B_n(n2693_n), .Y_n(n3395_n), .Y(n3395) );
 wddl_and U2220 ( .A(n2550), .A_n(n2550_n), .B(n2862), .B_n(n2862_n), .Y_n(n3394_n), .Y(n3394) );
 wddl_or U2221 ( .A(n2683), .A_n(n2683_n), .B(n2561), .B_n(n2561_n), .Y_n(n2862_n), .Y(n2862) );
 wddl_or U2222 ( .A(n3396), .A_n(n3396_n), .B(n3397), .B_n(n3397_n), .Y_n(n3392_n), .Y(n3392) );
 wddl_and U2223 ( .A(n2799), .A_n(n2799_n), .B(n2967), .B_n(n2967_n), .Y_n(n3397_n), .Y(n3397) );
 wddl_or U2224 ( .A(n2536), .A_n(n2536_n), .B(n2550), .B_n(n2550_n), .Y_n(n2967_n), .Y(n2967) );
 wddl_and U2225 ( .A(n2576), .A_n(n2576_n), .B(n2969), .B_n(n2969_n), .Y_n(n3396_n), .Y(n3396) );
 wddl_or U2226 ( .A(n2610), .A_n(n2610_n), .B(n2586), .B_n(n2586_n), .Y_n(n2969_n), .Y(n2969) );
 wddl_and U2227 ( .A(n2639), .A_n(n2639_n), .B(n3398), .B_n(n3398_n), .Y_n(n3390_n), .Y(n3390) );
 wddl_or U2228 ( .A(n2609), .A_n(n2609_n), .B(n3080), .B_n(n3080_n), .Y_n(n3398_n), .Y(n3398) );
 wddl_or U2229 ( .A(n3399), .A_n(n3399_n), .B(n3400), .B_n(n3400_n), .Y_n(n2851_n), .Y(n2851) );
 wddl_or U2230 ( .A(n3401), .A_n(n3401_n), .B(n3402), .B_n(n3402_n), .Y_n(n3400_n), .Y(n3400) );
 wddl_or U2231 ( .A(n3223), .A_n(n3223_n), .B(n3403), .B_n(n3403_n), .Y_n(n3402_n), .Y(n3402) );
 wddl_or U2232 ( .A(n3404), .A_n(n3404_n), .B(n3405), .B_n(n3405_n), .Y_n(n3403_n), .Y(n3403) );
 wddl_and U2233 ( .A(n2772), .A_n(n2772_n), .B(n2645), .B_n(n2645_n), .Y_n(n3405_n), .Y(n3405) );
 wddl_and U2234 ( .A(n2606), .A_n(n2606_n), .B(n2701), .B_n(n2701_n), .Y_n(n3404_n), .Y(n3404) );
 wddl_and U2235 ( .A(n2679), .A_n(n2679_n), .B(n2633), .B_n(n2633_n), .Y_n(n3401_n), .Y(n3401) );
 wddl_or U2236 ( .A(n3406), .A_n(n3406_n), .B(n3407), .B_n(n3407_n), .Y_n(n3399_n), .Y(n3399) );
 wddl_or U2237 ( .A(n3408), .A_n(n3408_n), .B(n3409), .B_n(n3409_n), .Y_n(n3407_n), .Y(n3407) );
 wddl_and U2238 ( .A(n2561), .A_n(n2561_n), .B(n2911), .B_n(n2911_n), .Y_n(n3409_n), .Y(n3409) );
 wddl_or U2239 ( .A(n2570), .A_n(n2570_n), .B(n3410), .B_n(n3410_n), .Y_n(n2911_n), .Y(n2911) );
 wddl_or U2240 ( .A(n2650), .A_n(n2650_n), .B(n2698), .B_n(n2698_n), .Y_n(n3410_n), .Y(n3410) );
 wddl_and U2241 ( .A(n2760), .A_n(n2760_n), .B(n3274), .B_n(n3274_n), .Y_n(n3408_n), .Y(n3408) );
 wddl_or U2242 ( .A(n3415), .A_n(n3415_n), .B(n3416), .B_n(n3416_n), .Y_n(n3406_n), .Y(n3406) );
 wddl_or U2243 ( .A(n3417), .A_n(n3417_n), .B(n3418), .B_n(n3418_n), .Y_n(n3416_n), .Y(n3416) );
 wddl_and U2244 ( .A(n2665), .A_n(n2665_n), .B(n3419), .B_n(n3419_n), .Y_n(n3418_n), .Y(n3418) );
 wddl_or U2245 ( .A(n2691), .A_n(n2691_n), .B(n2638), .B_n(n2638_n), .Y_n(n3419_n), .Y(n3419) );
 wddl_and U2246 ( .A(n2693), .A_n(n2693_n), .B(n3421), .B_n(n3421_n), .Y_n(n3417_n), .Y(n3417) );
 wddl_or U2247 ( .A(n2542), .A_n(n2542_n), .B(n2559), .B_n(n2559_n), .Y_n(n3421_n), .Y(n3421) );
 wddl_and U2248 ( .A(n2628), .A_n(n2628_n), .B(n3422), .B_n(n3422_n), .Y_n(n3415_n), .Y(n3415) );
 wddl_or U2249 ( .A(n2620), .A_n(n2620_n), .B(n2856), .B_n(n2856_n), .Y_n(n3422_n), .Y(n3422) );
 wddl_or U2250 ( .A(n2584), .A_n(n2584_n), .B(n2656), .B_n(n2656_n), .Y_n(n2856_n), .Y(n2856) );
 wddl_or U2251 ( .A(n3023), .A_n(n3023_n), .B(n3425), .B_n(n3425_n), .Y_n(n3362_n), .Y(n3362) );
 wddl_or U2252 ( .A(n3426), .A_n(n3426_n), .B(n3427), .B_n(n3427_n), .Y_n(n3425_n), .Y(n3425) );
 wddl_or U2253 ( .A(n3428), .A_n(n3428_n), .B(n3429), .B_n(n3429_n), .Y_n(n3427_n), .Y(n3427) );
 wddl_and U2254 ( .A(n2805), .A_n(n2805_n), .B(n2611), .B_n(n2611_n), .Y_n(n3429_n), .Y(n3429) );
 wddl_and U2255 ( .A(n2660), .A_n(n2660_n), .B(n2640), .B_n(n2640_n), .Y_n(n3428_n), .Y(n3428) );
 wddl_and U2256 ( .A(n2709), .A_n(n2709_n), .B(n3049), .B_n(n3049_n), .Y_n(n3426_n), .Y(n3426) );
 wddl_or U2257 ( .A(n3433), .A_n(n3433_n), .B(n3434), .B_n(n3434_n), .Y_n(n3023_n), .Y(n3023) );
 wddl_or U2258 ( .A(n3435), .A_n(n3435_n), .B(n3436), .B_n(n3436_n), .Y_n(n3434_n), .Y(n3434) );
 wddl_or U2259 ( .A(n3437), .A_n(n3437_n), .B(n3438), .B_n(n3438_n), .Y_n(n3436_n), .Y(n3436) );
 wddl_and U2260 ( .A(n2620), .A_n(n2620_n), .B(n2788), .B_n(n2788_n), .Y_n(n3438_n), .Y(n3438) );
 wddl_and U2261 ( .A(n2655), .A_n(n2655_n), .B(n2979), .B_n(n2979_n), .Y_n(n3437_n), .Y(n3437) );
 wddl_or U2262 ( .A(n2558), .A_n(n2558_n), .B(n2575), .B_n(n2575_n), .Y_n(n2979_n), .Y(n2979) );
 wddl_or U2263 ( .A(n3279), .A_n(n3279_n), .B(n3442), .B_n(n3442_n), .Y_n(n3435_n), .Y(n3435) );
 wddl_and U2264 ( .A(n2651), .A_n(n2651_n), .B(n3443), .B_n(n3443_n), .Y_n(n3442_n), .Y(n3442) );
 wddl_or U2265 ( .A(n2588), .A_n(n2588_n), .B(n2540), .B_n(n2540_n), .Y_n(n3443_n), .Y(n3443) );
 wddl_or U2266 ( .A(n3447), .A_n(n3447_n), .B(n3448), .B_n(n3448_n), .Y_n(n3433_n), .Y(n3433) );
 wddl_or U2267 ( .A(n3449), .A_n(n3449_n), .B(n3450), .B_n(n3450_n), .Y_n(n3448_n), .Y(n3448) );
 wddl_and U2268 ( .A(n2635), .A_n(n2635_n), .B(n3451), .B_n(n3451_n), .Y_n(n3450_n), .Y(n3450) );
 wddl_or U2269 ( .A(n2707), .A_n(n2707_n), .B(n2839), .B_n(n2839_n), .Y_n(n3451_n), .Y(n3451) );
 wddl_or U2270 ( .A(n2578), .A_n(n2578_n), .B(n2562), .B_n(n2562_n), .Y_n(n2839_n), .Y(n2839) );
 wddl_and U2271 ( .A(n2536), .A_n(n2536_n), .B(n3453), .B_n(n3453_n), .Y_n(n3449_n), .Y(n3449) );
 wddl_or U2272 ( .A(n2773), .A_n(n2773_n), .B(n2555), .B_n(n2555_n), .Y_n(n3453_n), .Y(n3453) );
 wddl_or U2273 ( .A(n3455), .A_n(n3455_n), .B(n3456), .B_n(n3456_n), .Y_n(n3447_n), .Y(n3447) );
 wddl_and U2274 ( .A(n2542), .A_n(n2542_n), .B(n3457), .B_n(n3457_n), .Y_n(n3456_n), .Y(n3456) );
 wddl_or U2275 ( .A(n2625), .A_n(n2625_n), .B(n2765), .B_n(n2765_n), .Y_n(n3457_n), .Y(n3457) );
 wddl_or U2276 ( .A(n2599), .A_n(n2599_n), .B(n2593), .B_n(n2593_n), .Y_n(n2765_n), .Y(n2765) );
 wddl_and U2277 ( .A(n2641), .A_n(n2641_n), .B(n3458), .B_n(n3458_n), .Y_n(n3455_n), .Y(n3455) );
 wddl_or U2278 ( .A(n2675), .A_n(n2675_n), .B(n2601), .B_n(n2601_n), .Y_n(n3458_n), .Y(n3458) );
 wddl_or U2279 ( .A(n2876), .A_n(n2876_n), .B(n3114), .B_n(n3114_n), .Y_n(d_n[1]), .Y(d[1]) );
 wddl_or U2280 ( .A(n3115), .A_n(n3115_n), .B(n3116), .B_n(n3116_n), .Y_n(n3114_n), .Y(n3114) );
 wddl_or U2281 ( .A(n3117), .A_n(n3117_n), .B(n3118), .B_n(n3118_n), .Y_n(n3116_n), .Y(n3116) );
 wddl_or U2282 ( .A(n2734), .A_n(n2734_n), .B(n2779), .B_n(n2779_n), .Y_n(n3118_n), .Y(n3118) );
 wddl_or U2283 ( .A(n3119), .A_n(n3119_n), .B(n3120), .B_n(n3120_n), .Y_n(n2779_n), .Y(n2779) );
 wddl_or U2284 ( .A(n3121), .A_n(n3121_n), .B(n3122), .B_n(n3122_n), .Y_n(n3120_n), .Y(n3120) );
 wddl_or U2285 ( .A(n3123), .A_n(n3123_n), .B(n3124), .B_n(n3124_n), .Y_n(n3122_n), .Y(n3122) );
 wddl_and U2286 ( .A(n2681), .A_n(n2681_n), .B(n2696), .B_n(n2696_n), .Y_n(n3124_n), .Y(n3124) );
 wddl_and U2287 ( .A(n2557), .A_n(n2557_n), .B(n2811), .B_n(n2811_n), .Y_n(n3123_n), .Y(n3123) );
 wddl_or U2288 ( .A(n3125), .A_n(n3125_n), .B(n3126), .B_n(n3126_n), .Y_n(n3121_n), .Y(n3121) );
 wddl_or U2289 ( .A(n2866), .A_n(n2866_n), .B(n3127), .B_n(n3127_n), .Y_n(n3126_n), .Y(n3126) );
 wddl_and U2290 ( .A(n2756), .A_n(n2756_n), .B(n2663), .B_n(n2663_n), .Y_n(n3127_n), .Y(n3127) );
 wddl_and U2291 ( .A(n2629), .A_n(n2629_n), .B(n2609), .B_n(n2609_n), .Y_n(n2866_n), .Y(n2866) );
 wddl_and U2292 ( .A(n2615), .A_n(n2615_n), .B(n2641), .B_n(n2641_n), .Y_n(n3125_n), .Y(n3125) );
 wddl_or U2293 ( .A(n3128), .A_n(n3128_n), .B(n3129), .B_n(n3129_n), .Y_n(n3119_n), .Y(n3119) );
 wddl_or U2294 ( .A(n3130), .A_n(n3130_n), .B(n3131), .B_n(n3131_n), .Y_n(n3129_n), .Y(n3129) );
 wddl_or U2295 ( .A(n3132), .A_n(n3132_n), .B(n3133), .B_n(n3133_n), .Y_n(n3131_n), .Y(n3131) );
 wddl_and U2296 ( .A(n2822), .A_n(n2822_n), .B(n2939), .B_n(n2939_n), .Y_n(n3133_n), .Y(n3133) );
 wddl_or U2297 ( .A(n2709), .A_n(n2709_n), .B(n2554), .B_n(n2554_n), .Y_n(n2939_n), .Y(n2939) );
 wddl_and U2298 ( .A(n2618), .A_n(n2618_n), .B(n3134), .B_n(n3134_n), .Y_n(n3132_n), .Y(n3132) );
 wddl_or U2299 ( .A(n2563), .A_n(n2563_n), .B(n2669), .B_n(n2669_n), .Y_n(n3134_n), .Y(n3134) );
 wddl_or U2300 ( .A(n3135), .A_n(n3135_n), .B(n3136), .B_n(n3136_n), .Y_n(n3130_n), .Y(n3130) );
 wddl_and U2301 ( .A(n2703), .A_n(n2703_n), .B(n3048), .B_n(n3048_n), .Y_n(n3136_n), .Y(n3136) );
 wddl_or U2302 ( .A(n2569), .A_n(n2569_n), .B(n2811), .B_n(n2811_n), .Y_n(n3048_n), .Y(n3048) );
 wddl_and U2303 ( .A(n2566), .A_n(n2566_n), .B(n3137), .B_n(n3137_n), .Y_n(n3135_n), .Y(n3135) );
 wddl_and U2304 ( .A(n2749), .A_n(n2749_n), .B(n3138), .B_n(n3138_n), .Y_n(n3128_n), .Y(n3128) );
 wddl_or U2305 ( .A(n2589), .A_n(n2589_n), .B(n2526), .B_n(n2526_n), .Y_n(n3138_n), .Y(n3138) );
 wddl_or U2306 ( .A(n3139), .A_n(n3139_n), .B(n3140), .B_n(n3140_n), .Y_n(n2734_n), .Y(n2734) );
 wddl_or U2307 ( .A(n3141), .A_n(n3141_n), .B(n3142), .B_n(n3142_n), .Y_n(n3140_n), .Y(n3140) );
 wddl_or U2308 ( .A(n3143), .A_n(n3143_n), .B(n3144), .B_n(n3144_n), .Y_n(n3142_n), .Y(n3142) );
 wddl_and U2309 ( .A(n2670), .A_n(n2670_n), .B(n2653), .B_n(n2653_n), .Y_n(n3144_n), .Y(n3144) );
 wddl_and U2310 ( .A(n2600), .A_n(n2600_n), .B(n3145), .B_n(n3145_n), .Y_n(n3143_n), .Y(n3143) );
 wddl_or U2311 ( .A(n3146), .A_n(n3146_n), .B(n3147), .B_n(n3147_n), .Y_n(n3141_n), .Y(n3141) );
 wddl_or U2312 ( .A(n3148), .A_n(n3148_n), .B(n3059), .B_n(n3059_n), .Y_n(n3147_n), .Y(n3147) );
 wddl_and U2313 ( .A(n2675), .A_n(n2675_n), .B(n2567), .B_n(n2567_n), .Y_n(n3059_n), .Y(n3059) );
 wddl_and U2314 ( .A(n2686), .A_n(n2686_n), .B(n3149), .B_n(n3149_n), .Y_n(n3148_n), .Y(n3148) );
 wddl_and U2315 ( .A(n2589), .A_n(n2589_n), .B(n2660), .B_n(n2660_n), .Y_n(n3146_n), .Y(n3146) );
 wddl_or U2316 ( .A(n3150), .A_n(n3150_n), .B(n3151), .B_n(n3151_n), .Y_n(n3139_n), .Y(n3139) );
 wddl_or U2317 ( .A(n3152), .A_n(n3152_n), .B(n3153), .B_n(n3153_n), .Y_n(n3151_n), .Y(n3151) );
 wddl_and U2318 ( .A(n2616), .A_n(n2616_n), .B(n2703), .B_n(n2703_n), .Y_n(n3153_n), .Y(n3153) );
 wddl_and U2319 ( .A(n2698), .A_n(n2698_n), .B(n2761), .B_n(n2761_n), .Y_n(n3152_n), .Y(n3152) );
 wddl_or U2320 ( .A(n3154), .A_n(n3154_n), .B(n3155), .B_n(n3155_n), .Y_n(n3150_n), .Y(n3150) );
 wddl_or U2321 ( .A(n3156), .A_n(n3156_n), .B(n3157), .B_n(n3157_n), .Y_n(n3155_n), .Y(n3155) );
 wddl_and U2322 ( .A(n2688), .A_n(n2688_n), .B(n3158), .B_n(n3158_n), .Y_n(n3157_n), .Y(n3157) );
 wddl_or U2323 ( .A(n2674), .A_n(n2674_n), .B(n2569), .B_n(n2569_n), .Y_n(n3158_n), .Y(n3158) );
 wddl_and U2324 ( .A(n2575), .A_n(n2575_n), .B(n2800), .B_n(n2800_n), .Y_n(n3156_n), .Y(n3156) );
 wddl_or U2325 ( .A(n2538), .A_n(n2538_n), .B(n2659), .B_n(n2659_n), .Y_n(n2800_n), .Y(n2800) );
 wddl_and U2326 ( .A(n2635), .A_n(n2635_n), .B(n2745), .B_n(n2745_n), .Y_n(n3154_n), .Y(n3154) );
 wddl_and U2327 ( .A(n3159), .A_n(n3159_n), .B(n2715), .B_n(n2715_n), .Y_n(n2745_n), .Y(n2745) );
 wddl_or U2328 ( .A(n3160), .A_n(n3160_n), .B(n3161), .B_n(n3161_n), .Y_n(n3117_n), .Y(n3117) );
 wddl_or U2329 ( .A(n3162), .A_n(n3162_n), .B(n3163), .B_n(n3163_n), .Y_n(n3161_n), .Y(n3161) );
 wddl_and U2330 ( .A(n2629), .A_n(n2629_n), .B(n3164), .B_n(n3164_n), .Y_n(n3163_n), .Y(n3163) );
 wddl_or U2331 ( .A(n2594), .A_n(n2594_n), .B(n3080), .B_n(n3080_n), .Y_n(n3164_n), .Y(n3164) );
 wddl_or U2332 ( .A(n2626), .A_n(n2626_n), .B(n2636), .B_n(n2636_n), .Y_n(n3080_n), .Y(n3080) );
 wddl_and U2333 ( .A(n2645), .A_n(n2645_n), .B(n3165), .B_n(n3165_n), .Y_n(n3162_n), .Y(n3162) );
 wddl_or U2334 ( .A(n2648), .A_n(n2648_n), .B(n2664), .B_n(n2664_n), .Y_n(n3165_n), .Y(n3165) );
 wddl_or U2335 ( .A(n3166), .A_n(n3166_n), .B(n3167), .B_n(n3167_n), .Y_n(n3160_n), .Y(n3160) );
 wddl_or U2336 ( .A(n3168), .A_n(n3168_n), .B(n3169), .B_n(n3169_n), .Y_n(n3167_n), .Y(n3167) );
 wddl_or U2337 ( .A(n3170), .A_n(n3170_n), .B(n3171), .B_n(n3171_n), .Y_n(n3169_n), .Y(n3169) );
 wddl_or U2338 ( .A(n3172), .A_n(n3172_n), .B(n3173), .B_n(n3173_n), .Y_n(n3171_n), .Y(n3171) );
 wddl_and U2339 ( .A(n2559), .A_n(n2559_n), .B(n2585), .B_n(n2585_n), .Y_n(n3173_n), .Y(n3173) );
 wddl_and U2340 ( .A(n2685), .A_n(n2685_n), .B(n2570), .B_n(n2570_n), .Y_n(n3172_n), .Y(n3172) );
 wddl_and U2341 ( .A(n2573), .A_n(n2573_n), .B(n2655), .B_n(n2655_n), .Y_n(n3170_n), .Y(n3170) );
 wddl_and U2342 ( .A(n2688), .A_n(n2688_n), .B(n2836), .B_n(n2836_n), .Y_n(n3168_n), .Y(n3168) );
 wddl_or U2343 ( .A(n2613), .A_n(n2613_n), .B(n2583), .B_n(n2583_n), .Y_n(n2836_n), .Y(n2836) );
 wddl_and U2344 ( .A(n2615), .A_n(n2615_n), .B(n3174), .B_n(n3174_n), .Y_n(n3166_n), .Y(n3166) );
 wddl_or U2345 ( .A(n2588), .A_n(n2588_n), .B(n2888), .B_n(n2888_n), .Y_n(n3174_n), .Y(n3174) );
 wddl_or U2346 ( .A(n2645), .A_n(n2645_n), .B(n2678), .B_n(n2678_n), .Y_n(n2888_n), .Y(n2888) );
 wddl_or U2347 ( .A(n2843), .A_n(n2843_n), .B(n3175), .B_n(n3175_n), .Y_n(n3115_n), .Y(n3115) );
 wddl_or U2348 ( .A(n3051), .A_n(n3051_n), .B(n3176), .B_n(n3176_n), .Y_n(n3175_n), .Y(n3175) );
 wddl_or U2349 ( .A(n3177), .A_n(n3177_n), .B(n3178), .B_n(n3178_n), .Y_n(n3176_n), .Y(n3176) );
 wddl_and U2350 ( .A(n2611), .A_n(n2611_n), .B(n2639), .B_n(n2639_n), .Y_n(n3178_n), .Y(n3178) );
 wddl_and U2351 ( .A(n2565), .A_n(n2565_n), .B(n2658), .B_n(n2658_n), .Y_n(n3177_n), .Y(n3177) );
 wddl_and U2352 ( .A(n2708), .A_n(n2708_n), .B(n2623), .B_n(n2623_n), .Y_n(n3051_n), .Y(n3051) );
 wddl_or U2353 ( .A(n3179), .A_n(n3179_n), .B(n3180), .B_n(n3180_n), .Y_n(n2843_n), .Y(n2843) );
 wddl_or U2354 ( .A(n3181), .A_n(n3181_n), .B(n3182), .B_n(n3182_n), .Y_n(n3180_n), .Y(n3180) );
 wddl_or U2355 ( .A(n3183), .A_n(n3183_n), .B(n3095), .B_n(n3095_n), .Y_n(n3182_n), .Y(n3182) );
 wddl_and U2356 ( .A(n2624), .A_n(n2624_n), .B(n2588), .B_n(n2588_n), .Y_n(n3095_n), .Y(n3095) );
 wddl_and U2357 ( .A(n2741), .A_n(n2741_n), .B(n2584), .B_n(n2584_n), .Y_n(n3183_n), .Y(n3183) );
 wddl_or U2358 ( .A(n3184), .A_n(n3184_n), .B(n3185), .B_n(n3185_n), .Y_n(n3181_n), .Y(n3181) );
 wddl_and U2359 ( .A(n2634), .A_n(n2634_n), .B(n3145), .B_n(n3145_n), .Y_n(n3185_n), .Y(n3185) );
 wddl_or U2360 ( .A(n2580), .A_n(n2580_n), .B(n2557), .B_n(n2557_n), .Y_n(n3145_n), .Y(n3145) );
 wddl_and U2361 ( .A(n2613), .A_n(n2613_n), .B(n2575), .B_n(n2575_n), .Y_n(n3184_n), .Y(n3184) );
 wddl_or U2362 ( .A(n3186), .A_n(n3186_n), .B(n3187), .B_n(n3187_n), .Y_n(n3179_n), .Y(n3179) );
 wddl_or U2363 ( .A(n3188), .A_n(n3188_n), .B(n3189), .B_n(n3189_n), .Y_n(n3187_n), .Y(n3187) );
 wddl_and U2364 ( .A(n2595), .A_n(n2595_n), .B(n3190), .B_n(n3190_n), .Y_n(n3189_n), .Y(n3189) );
 wddl_or U2365 ( .A(n2681), .A_n(n2681_n), .B(n3191), .B_n(n3191_n), .Y_n(n3190_n), .Y(n3190) );
 wddl_or U2366 ( .A(n2703), .A_n(n2703_n), .B(n2771), .B_n(n2771_n), .Y_n(n3191_n), .Y(n3191) );
 wddl_and U2367 ( .A(n2559), .A_n(n2559_n), .B(n3192), .B_n(n3192_n), .Y_n(n3188_n), .Y(n3188) );
 wddl_or U2368 ( .A(n2701), .A_n(n2701_n), .B(n3137), .B_n(n3137_n), .Y_n(n3192_n), .Y(n3192) );
 wddl_or U2369 ( .A(n2693), .A_n(n2693_n), .B(n2874), .B_n(n2874_n), .Y_n(n3137_n), .Y(n3137) );
 wddl_or U2370 ( .A(n3193), .A_n(n3193_n), .B(n3194), .B_n(n3194_n), .Y_n(n3186_n), .Y(n3186) );
 wddl_and U2371 ( .A(n2683), .A_n(n2683_n), .B(n3195), .B_n(n3195_n), .Y_n(n3194_n), .Y(n3194) );
 wddl_or U2372 ( .A(n2651), .A_n(n2651_n), .B(n2990), .B_n(n2990_n), .Y_n(n3195_n), .Y(n3195) );
 wddl_or U2373 ( .A(n2635), .A_n(n2635_n), .B(n2829), .B_n(n2829_n), .Y_n(n2990_n), .Y(n2990) );
 wddl_and U2374 ( .A(n2546), .A_n(n2546_n), .B(n3196), .B_n(n3196_n), .Y_n(n3193_n), .Y(n3193) );
 wddl_or U2375 ( .A(n2555), .A_n(n2555_n), .B(n2563), .B_n(n2563_n), .Y_n(n3196_n), .Y(n3196) );
 wddl_or U2376 ( .A(n3197), .A_n(n3197_n), .B(n3198), .B_n(n3198_n), .Y_n(n2876_n), .Y(n2876) );
 wddl_or U2377 ( .A(n2777), .A_n(n2777_n), .B(n3199), .B_n(n3199_n), .Y_n(n3198_n), .Y(n3198) );
 wddl_or U2378 ( .A(n2816), .A_n(n2816_n), .B(n3200), .B_n(n3200_n), .Y_n(n3199_n), .Y(n3199) );
 wddl_or U2379 ( .A(n3201), .A_n(n3201_n), .B(n3202), .B_n(n3202_n), .Y_n(n3200_n), .Y(n3200) );
 wddl_or U2380 ( .A(n3203), .A_n(n3203_n), .B(n3204), .B_n(n3204_n), .Y_n(n3202_n), .Y(n3202) );
 wddl_or U2381 ( .A(n3205), .A_n(n3205_n), .B(n3206), .B_n(n3206_n), .Y_n(n3204_n), .Y(n3204) );
 wddl_and U2382 ( .A(n2648), .A_n(n2648_n), .B(n2746), .B_n(n2746_n), .Y_n(n3206_n), .Y(n3206) );
 wddl_and U2383 ( .A(n2524), .A_n(n2524_n), .B(n3299), .B_n(n3299_n), .Y_n(n2746_n), .Y(n2746) );
 wddl_and U2384 ( .A(n2710), .A_n(n2710_n), .B(n2636), .B_n(n2636_n), .Y_n(n3205_n), .Y(n3205) );
 wddl_and U2385 ( .A(n2625), .A_n(n2625_n), .B(n2563), .B_n(n2563_n), .Y_n(n3203_n), .Y(n3203) );
 wddl_and U2386 ( .A(n2533), .A_n(n2533_n), .B(n2531), .B_n(n2531_n), .Y_n(n2770_n), .Y(n2770) );
 wddl_or U2387 ( .A(n3207), .A_n(n3207_n), .B(n3208), .B_n(n3208_n), .Y_n(n3201_n), .Y(n3201) );
 wddl_or U2388 ( .A(n3209), .A_n(n3209_n), .B(n3210), .B_n(n3210_n), .Y_n(n3208_n), .Y(n3208) );
 wddl_or U2389 ( .A(n3211), .A_n(n3211_n), .B(n3212), .B_n(n3212_n), .Y_n(n3210_n), .Y(n3210) );
 wddl_and U2390 ( .A(n2631), .A_n(n2631_n), .B(n3213), .B_n(n3213_n), .Y_n(n3212_n), .Y(n3212) );
 wddl_or U2391 ( .A(n2696), .A_n(n2696_n), .B(n2665), .B_n(n2665_n), .Y_n(n3213_n), .Y(n3213) );
 wddl_and U2392 ( .A(n2690), .A_n(n2690_n), .B(n3214), .B_n(n3214_n), .Y_n(n3211_n), .Y(n3211) );
 wddl_or U2393 ( .A(n2598), .A_n(n2598_n), .B(n2699), .B_n(n2699_n), .Y_n(n3214_n), .Y(n3214) );
 wddl_and U2394 ( .A(n2571), .A_n(n2571_n), .B(n3215), .B_n(n3215_n), .Y_n(n3209_n), .Y(n3209) );
 wddl_or U2395 ( .A(n2799), .A_n(n2799_n), .B(n2573), .B_n(n2573_n), .Y_n(n3215_n), .Y(n3215) );
 wddl_and U2396 ( .A(n2614), .A_n(n2614_n), .B(n3216), .B_n(n3216_n), .Y_n(n3207_n), .Y(n3207) );
 wddl_or U2397 ( .A(n2603), .A_n(n2603_n), .B(n2671), .B_n(n2671_n), .Y_n(n3216_n), .Y(n3216) );
 wddl_or U2398 ( .A(n3217), .A_n(n3217_n), .B(n3218), .B_n(n3218_n), .Y_n(n2816_n), .Y(n2816) );
 wddl_or U2399 ( .A(n3219), .A_n(n3219_n), .B(n3220), .B_n(n3220_n), .Y_n(n3218_n), .Y(n3218) );
 wddl_or U2400 ( .A(n3221), .A_n(n3221_n), .B(n3222), .B_n(n3222_n), .Y_n(n3220_n), .Y(n3220) );
 wddl_or U2401 ( .A(n3223), .A_n(n3223_n), .B(n3224), .B_n(n3224_n), .Y_n(n3222_n), .Y(n3222) );
 wddl_and U2402 ( .A(n2567), .A_n(n2567_n), .B(n2701), .B_n(n2701_n), .Y_n(n3224_n), .Y(n3224) );
 wddl_and U2403 ( .A(n2570), .A_n(n2570_n), .B(n2548), .B_n(n2548_n), .Y_n(n3223_n), .Y(n3223) );
 wddl_and U2404 ( .A(n2610), .A_n(n2610_n), .B(n2761), .B_n(n2761_n), .Y_n(n3221_n), .Y(n3221) );
 wddl_or U2405 ( .A(n2562), .A_n(n2562_n), .B(n2576), .B_n(n2576_n), .Y_n(n2761_n), .Y(n2761) );
 wddl_and U2406 ( .A(n2678), .A_n(n2678_n), .B(n2665), .B_n(n2665_n), .Y_n(n3219_n), .Y(n3219) );
 wddl_or U2407 ( .A(n3225), .A_n(n3225_n), .B(n3226), .B_n(n3226_n), .Y_n(n3217_n), .Y(n3217) );
 wddl_or U2408 ( .A(n3227), .A_n(n3227_n), .B(n3228), .B_n(n3228_n), .Y_n(n3226_n), .Y(n3226) );
 wddl_and U2409 ( .A(n2649), .A_n(n2649_n), .B(n2522), .B_n(n2522_n), .Y_n(n3228_n), .Y(n3228) );
 wddl_and U2410 ( .A(n2586), .A_n(n2586_n), .B(n3229), .B_n(n3229_n), .Y_n(n3227_n), .Y(n3227) );
 wddl_or U2411 ( .A(n2678), .A_n(n2678_n), .B(n2640), .B_n(n2640_n), .Y_n(n3229_n), .Y(n3229) );
 wddl_or U2412 ( .A(n3230), .A_n(n3230_n), .B(n3231), .B_n(n3231_n), .Y_n(n3225_n), .Y(n3225) );
 wddl_or U2413 ( .A(n3232), .A_n(n3232_n), .B(n3233), .B_n(n3233_n), .Y_n(n3231_n), .Y(n3231) );
 wddl_and U2414 ( .A(n2646), .A_n(n2646_n), .B(n3234), .B_n(n3234_n), .Y_n(n3233_n), .Y(n3233) );
 wddl_or U2415 ( .A(n2619), .A_n(n2619_n), .B(n2658), .B_n(n2658_n), .Y_n(n3234_n), .Y(n3234) );
 wddl_and U2416 ( .A(n2709), .A_n(n2709_n), .B(n3235), .B_n(n3235_n), .Y_n(n3232_n), .Y(n3232) );
 wddl_or U2417 ( .A(n3149), .A_n(n3149_n), .B(n2618), .B_n(n2618_n), .Y_n(n3235_n), .Y(n3235) );
 wddl_and U2418 ( .A(n2691), .A_n(n2691_n), .B(n3236), .B_n(n3236_n), .Y_n(n3230_n), .Y(n3230) );
 wddl_or U2419 ( .A(n2634), .A_n(n2634_n), .B(n2655), .B_n(n2655_n), .Y_n(n3236_n), .Y(n3236) );
 wddl_or U2420 ( .A(n3237), .A_n(n3237_n), .B(n3238), .B_n(n3238_n), .Y_n(n2777_n), .Y(n2777) );
 wddl_or U2421 ( .A(n3239), .A_n(n3239_n), .B(n3240), .B_n(n3240_n), .Y_n(n3238_n), .Y(n3238) );
 wddl_or U2422 ( .A(n3241), .A_n(n3241_n), .B(n3242), .B_n(n3242_n), .Y_n(n3240_n), .Y(n3240) );
 wddl_and U2423 ( .A(n2593), .A_n(n2593_n), .B(n2669), .B_n(n2669_n), .Y_n(n3242_n), .Y(n3242) );
 wddl_and U2424 ( .A(n2650), .A_n(n2650_n), .B(n2690), .B_n(n2690_n), .Y_n(n3241_n), .Y(n3241) );
 wddl_or U2425 ( .A(n3243), .A_n(n3243_n), .B(n3244), .B_n(n3244_n), .Y_n(n3239_n), .Y(n3239) );
 wddl_and U2426 ( .A(n2707), .A_n(n2707_n), .B(n2666), .B_n(n2666_n), .Y_n(n3244_n), .Y(n3244) );
 wddl_and U2427 ( .A(n2895), .A_n(n2895_n), .B(n3112), .B_n(n3112_n), .Y_n(n3243_n), .Y(n3243) );
 wddl_or U2428 ( .A(n2646), .A_n(n2646_n), .B(n2669), .B_n(n2669_n), .Y_n(n3112_n), .Y(n3112) );
 wddl_and U2429 ( .A(n3439), .A_n(n3439_n), .B(n3413), .B_n(n3413_n), .Y_n(n2788_n), .Y(n2788) );
 wddl_or U2430 ( .A(n3245), .A_n(n3245_n), .B(n3246), .B_n(n3246_n), .Y_n(n3237_n), .Y(n3237) );
 wddl_or U2431 ( .A(n3247), .A_n(n3247_n), .B(n3248), .B_n(n3248_n), .Y_n(n3246_n), .Y(n3246) );
 wddl_and U2432 ( .A(n2600), .A_n(n2600_n), .B(n3249), .B_n(n3249_n), .Y_n(n3248_n), .Y(n3248) );
 wddl_or U2433 ( .A(n2630), .A_n(n2630_n), .B(n2544), .B_n(n2544_n), .Y_n(n3249_n), .Y(n3249) );
 wddl_and U2434 ( .A(n3452), .A_n(n3452_n), .B(n3440), .B_n(n3440_n), .Y_n(n2822_n), .Y(n2822) );
 wddl_and U2435 ( .A(n2608), .A_n(n2608_n), .B(n2863), .B_n(n2863_n), .Y_n(n3247_n), .Y(n3247) );
 wddl_and U2436 ( .A(n2524), .A_n(n2524_n), .B(n3251), .B_n(n3251_n), .Y_n(n2863_n), .Y(n2863) );
 wddl_or U2437 ( .A(n3252), .A_n(n3252_n), .B(n3253), .B_n(n3253_n), .Y_n(n3245_n), .Y(n3245) );
 wddl_or U2438 ( .A(n3254), .A_n(n3254_n), .B(n3255), .B_n(n3255_n), .Y_n(n3253_n), .Y(n3253) );
 wddl_and U2439 ( .A(n2659), .A_n(n2659_n), .B(n3256), .B_n(n3256_n), .Y_n(n3255_n), .Y(n3255) );
 wddl_or U2440 ( .A(n2629), .A_n(n2629_n), .B(n2797), .B_n(n2797_n), .Y_n(n3256_n), .Y(n3256) );
 wddl_and U2441 ( .A(n3430), .A_n(n3430_n), .B(n3431), .B_n(n3431_n), .Y_n(n2811_n), .Y(n2811) );
 wddl_and U2442 ( .A(n2723), .A_n(n2723_n), .B(n3424), .B_n(n3424_n), .Y_n(n3431_n), .Y(n3431) );
 wddl_and U2443 ( .A(n2653), .A_n(n2653_n), .B(n3257), .B_n(n3257_n), .Y_n(n3254_n), .Y(n3254) );
 wddl_or U2444 ( .A(n2580), .A_n(n2580_n), .B(n2565), .B_n(n2565_n), .Y_n(n3257_n), .Y(n3257) );
 wddl_and U2445 ( .A(n2621), .A_n(n2621_n), .B(n3258), .B_n(n3258_n), .Y_n(n3252_n), .Y(n3252) );
 wddl_or U2446 ( .A(n2574), .A_n(n2574_n), .B(n2897), .B_n(n2897_n), .Y_n(n3258_n), .Y(n3258) );
 wddl_or U2447 ( .A(n2631), .A_n(n2631_n), .B(n2603), .B_n(n2603_n), .Y_n(n2897_n), .Y(n2897) );
 wddl_or U2448 ( .A(n2766), .A_n(n2766_n), .B(n3259), .B_n(n3259_n), .Y_n(n3197_n), .Y(n3197) );
 wddl_or U2449 ( .A(n3260), .A_n(n3260_n), .B(n3261), .B_n(n3261_n), .Y_n(n3259_n), .Y(n3259) );
 wddl_or U2450 ( .A(n3262), .A_n(n3262_n), .B(n3263), .B_n(n3263_n), .Y_n(n3261_n), .Y(n3261) );
 wddl_or U2451 ( .A(n3264), .A_n(n3264_n), .B(n3265), .B_n(n3265_n), .Y_n(n3263_n), .Y(n3263) );
 wddl_and U2452 ( .A(n2686), .A_n(n2686_n), .B(n2694), .B_n(n2694_n), .Y_n(n3265_n), .Y(n3265) );
 wddl_and U2453 ( .A(n3444), .A_n(n3444_n), .B(n2524), .B_n(n2524_n), .Y_n(n2756_n), .Y(n2756) );
 wddl_and U2454 ( .A(n2554), .A_n(n2554_n), .B(n2619), .B_n(n2619_n), .Y_n(n3264_n), .Y(n3264) );
 wddl_and U2455 ( .A(n3440), .A_n(n3440_n), .B(n3412), .B_n(n3412_n), .Y_n(n2874_n), .Y(n2874) );
 wddl_and U2456 ( .A(n3414), .A_n(n3414_n), .B(n3441), .B_n(n3441_n), .Y_n(n2805_n), .Y(n2805) );
 wddl_and U2457 ( .A(n2581), .A_n(n2581_n), .B(n3049), .B_n(n3049_n), .Y_n(n3262_n), .Y(n3262) );
 wddl_or U2458 ( .A(n2593), .A_n(n2593_n), .B(n2611), .B_n(n2611_n), .Y_n(n3049_n), .Y(n3049) );
 wddl_and U2459 ( .A(n2681), .A_n(n2681_n), .B(n2610), .B_n(n2610_n), .Y_n(n3260_n), .Y(n3260) );
 wddl_and U2460 ( .A(n3430), .A_n(n3430_n), .B(n3432), .B_n(n3432_n), .Y_n(n2829_n), .Y(n2829) );
 wddl_and U2461 ( .A(n2726), .A_n(n2726_n), .B(n2724), .B_n(n2724_n), .Y_n(n3432_n), .Y(n3432) );
 wddl_or U2462 ( .A(n3266), .A_n(n3266_n), .B(n3267), .B_n(n3267_n), .Y_n(n2766_n), .Y(n2766) );
 wddl_or U2463 ( .A(n3268), .A_n(n3268_n), .B(n3269), .B_n(n3269_n), .Y_n(n3267_n), .Y(n3267) );
 wddl_or U2464 ( .A(n3270), .A_n(n3270_n), .B(n3271), .B_n(n3271_n), .Y_n(n3269_n), .Y(n3269) );
 wddl_and U2465 ( .A(n2678), .A_n(n2678_n), .B(n3065), .B_n(n3065_n), .Y_n(n3271_n), .Y(n3271) );
 wddl_or U2466 ( .A(n2546), .A_n(n2546_n), .B(n2536), .B_n(n2536_n), .Y_n(n3065_n), .Y(n3065) );
 wddl_and U2467 ( .A(n3430), .A_n(n3430_n), .B(n3454), .B_n(n3454_n), .Y_n(n2895_n), .Y(n2895) );
 wddl_and U2468 ( .A(n2534), .A_n(n2534_n), .B(n3380), .B_n(n3380_n), .Y_n(n3454_n), .Y(n3454) );
 wddl_and U2469 ( .A(n2718), .A_n(n2718_n), .B(n2995), .B_n(n2995_n), .Y_n(n2804_n), .Y(n2804) );
 wddl_and U2470 ( .A(n2580), .A_n(n2580_n), .B(n3085), .B_n(n3085_n), .Y_n(n3270_n), .Y(n3270) );
 wddl_or U2471 ( .A(n2676), .A_n(n2676_n), .B(n2666), .B_n(n2666_n), .Y_n(n3085_n), .Y(n3085) );
 wddl_and U2472 ( .A(n3412), .A_n(n3412_n), .B(n3420), .B_n(n3420_n), .Y_n(n2786_n), .Y(n2786) );
 wddl_and U2473 ( .A(n2722), .A_n(n2722_n), .B(n2723), .B_n(n2723_n), .Y_n(n3420_n), .Y(n3420) );
 wddl_and U2474 ( .A(n3430), .A_n(n3430_n), .B(n3459), .B_n(n3459_n), .Y_n(n2772_n), .Y(n2772) );
 wddl_and U2475 ( .A(n2531), .A_n(n2531_n), .B(n2725), .B_n(n2725_n), .Y_n(n3459_n), .Y(n3459) );
 wddl_and U2476 ( .A(n2722), .A_n(n2722_n), .B(n2720), .B_n(n2720_n), .Y_n(n3430_n), .Y(n3430) );
 wddl_and U2477 ( .A(n3441), .A_n(n3441_n), .B(n2528), .B_n(n2528_n), .Y_n(n2798_n), .Y(n2798) );
 wddl_or U2478 ( .A(n3272), .A_n(n3272_n), .B(n3273), .B_n(n3273_n), .Y_n(n3268_n), .Y(n3268) );
 wddl_and U2479 ( .A(n3439), .A_n(n3439_n), .B(n3414), .B_n(n3414_n), .Y_n(n2799_n), .Y(n2799) );
 wddl_and U2480 ( .A(n2758), .A_n(n2758_n), .B(n3380), .B_n(n3380_n), .Y_n(n2748_n), .Y(n2748) );
 wddl_and U2481 ( .A(n2722), .A_n(n2722_n), .B(n3452), .B_n(n3452_n), .Y_n(n2758_n), .Y(n2758) );
 wddl_and U2482 ( .A(n2636), .A_n(n2636_n), .B(n3274), .B_n(n3274_n), .Y_n(n3272_n), .Y(n3272) );
 wddl_or U2483 ( .A(n2643), .A_n(n2643_n), .B(n2567), .B_n(n2567_n), .Y_n(n3274_n), .Y(n3274) );
 wddl_and U2484 ( .A(n3250), .A_n(n3250_n), .B(n3414), .B_n(n3414_n), .Y_n(n2741_n), .Y(n2741) );
 wddl_and U2485 ( .A(n2716), .A_n(n2716_n), .B(n3251), .B_n(n3251_n), .Y_n(n3414_n), .Y(n3414) );
 wddl_and U2486 ( .A(n3452), .A_n(n3452_n), .B(n3411), .B_n(n3411_n), .Y_n(n2764_n), .Y(n2764) );
 wddl_and U2487 ( .A(n2726), .A_n(n2726_n), .B(n2719), .B_n(n2719_n), .Y_n(n3452_n), .Y(n3452) );
 wddl_or U2488 ( .A(n3275), .A_n(n3275_n), .B(n3276), .B_n(n3276_n), .Y_n(n3266_n), .Y(n3266) );
 wddl_or U2489 ( .A(n3277), .A_n(n3277_n), .B(n3278), .B_n(n3278_n), .Y_n(n3276_n), .Y(n3276) );
 wddl_or U2490 ( .A(n3279), .A_n(n3279_n), .B(n3280), .B_n(n3280_n), .Y_n(n3278_n), .Y(n3278) );
 wddl_and U2491 ( .A(n2655), .A_n(n2655_n), .B(n2638), .B_n(n2638_n), .Y_n(n3280_n), .Y(n3280) );
 wddl_and U2492 ( .A(n3444), .A_n(n3444_n), .B(n3159), .B_n(n3159_n), .Y_n(n2797_n), .Y(n2797) );
 wddl_and U2493 ( .A(n3149), .A_n(n3149_n), .B(n3424), .B_n(n3424_n), .Y_n(n2749_n), .Y(n2749) );
 wddl_and U2494 ( .A(n2590), .A_n(n2590_n), .B(n2695), .B_n(n2695_n), .Y_n(n3279_n), .Y(n3279) );
 wddl_and U2495 ( .A(n3412), .A_n(n3412_n), .B(n3446), .B_n(n3446_n), .Y_n(n2744_n), .Y(n2744) );
 wddl_and U2496 ( .A(n2722), .A_n(n2722_n), .B(n2724), .B_n(n2724_n), .Y_n(n3446_n), .Y(n3446) );
 wddl_or U2497 ( .A(n3281), .A_n(n3281_n), .B(n3282), .B_n(n3282_n), .Y_n(n3277_n), .Y(n3277) );
 wddl_or U2498 ( .A(n3283), .A_n(n3283_n), .B(n3097), .B_n(n3097_n), .Y_n(n3282_n), .Y(n3282) );
 wddl_and U2499 ( .A(n2760), .A_n(n2760_n), .B(n2605), .B_n(n2605_n), .Y_n(n3097_n), .Y(n3097) );
 wddl_and U2500 ( .A(n2528), .A_n(n2528_n), .B(n3159), .B_n(n3159_n), .Y_n(n2771_n), .Y(n2771) );
 wddl_and U2501 ( .A(n3411), .A_n(n3411_n), .B(n3445), .B_n(n3445_n), .Y_n(n2760_n), .Y(n2760) );
 wddl_and U2502 ( .A(n2534), .A_n(n2534_n), .B(n2720), .B_n(n2720_n), .Y_n(n3445_n), .Y(n3445) );
 wddl_and U2503 ( .A(n2583), .A_n(n2583_n), .B(n2530), .B_n(n2530_n), .Y_n(n3283_n), .Y(n3283) );
 wddl_or U2504 ( .A(n2567), .A_n(n2567_n), .B(n2573), .B_n(n2573_n), .Y_n(n2875_n), .Y(n2875) );
 wddl_and U2505 ( .A(n3441), .A_n(n3441_n), .B(n3413), .B_n(n3413_n), .Y_n(n2762_n), .Y(n2762) );
 wddl_and U2506 ( .A(n3250), .A_n(n3250_n), .B(n3413), .B_n(n3413_n), .Y_n(n2759_n), .Y(n2759) );
 wddl_and U2507 ( .A(n2718), .A_n(n2718_n), .B(n2716), .B_n(n2716_n), .Y_n(n3413_n), .Y(n3413) );
 wddl_and U2508 ( .A(n2712), .A_n(n2712_n), .B(n2713), .B_n(n2713_n), .Y_n(n3250_n), .Y(n3250) );
 wddl_and U2509 ( .A(n3411), .A_n(n3411_n), .B(n3423), .B_n(n3423_n), .Y_n(n2757_n), .Y(n2757) );
 wddl_and U2510 ( .A(n2720), .A_n(n2720_n), .B(n3424), .B_n(n3424_n), .Y_n(n3423_n), .Y(n3423) );
 wddl_and U2511 ( .A(n2596), .A_n(n2596_n), .B(n2830), .B_n(n2830_n), .Y_n(n3281_n), .Y(n3281) );
 wddl_and U2512 ( .A(n3444), .A_n(n3444_n), .B(n3441), .B_n(n3441_n), .Y_n(n2830_n), .Y(n2830) );
 wddl_and U2513 ( .A(n2714), .A_n(n2714_n), .B(n2711), .B_n(n2711_n), .Y_n(n3441_n), .Y(n3441) );
 wddl_and U2514 ( .A(n2726), .A_n(n2726_n), .B(n3149), .B_n(n3149_n), .Y_n(n2743_n), .Y(n2743) );
 wddl_and U2515 ( .A(n2720), .A_n(n2720_n), .B(n3440), .B_n(n3440_n), .Y_n(n3149_n), .Y(n3149) );
 wddl_and U2516 ( .A(n3380), .A_n(n3380_n), .B(n2721), .B_n(n2721_n), .Y_n(n3440_n), .Y(n3440) );
 wddl_and U2517 ( .A(n2796), .A_n(n2796_n), .B(n3284), .B_n(n3284_n), .Y_n(n3275_n), .Y(n3275) );
 wddl_or U2518 ( .A(n2629), .A_n(n2629_n), .B(n2900), .B_n(n2900_n), .Y_n(n3284_n), .Y(n3284) );
 wddl_or U2519 ( .A(n2589), .A_n(n2589_n), .B(n2561), .B_n(n2561_n), .Y_n(n2900_n), .Y(n2900) );
 wddl_and U2520 ( .A(n3439), .A_n(n3439_n), .B(n3299), .B_n(n3299_n), .Y_n(n2835_n), .Y(n2835) );
 wddl_and U2521 ( .A(n2715), .A_n(n2715_n), .B(n3251), .B_n(n3251_n), .Y_n(n3299_n), .Y(n3299) );
 wddl_and U2522 ( .A(n2522), .A_n(n2522_n), .B(n3251), .B_n(n3251_n), .Y_n(n2868_n), .Y(n2868) );
 wddl_and U2523 ( .A(n2716), .A_n(n2716_n), .B(n3159), .B_n(n3159_n), .Y_n(n2995_n), .Y(n2995) );
 wddl_and U2524 ( .A(n2712), .A_n(n2712_n), .B(n2714), .B_n(n2714_n), .Y_n(n3159_n), .Y(n3159) );
 wddl_and U2525 ( .A(n3444), .A_n(n3444_n), .B(n3439), .B_n(n3439_n), .Y_n(n2773_n), .Y(n2773) );
 wddl_and U2526 ( .A(n2713), .A_n(n2713_n), .B(n2711), .B_n(n2711_n), .Y_n(n3439_n), .Y(n3439) );
 wddl_and U2527 ( .A(n2718), .A_n(n2718_n), .B(n2715), .B_n(n2715_n), .Y_n(n3444_n), .Y(n3444) );
 wddl_and U2528 ( .A(n3411), .A_n(n3411_n), .B(n3412), .B_n(n3412_n), .Y_n(n2796_n), .Y(n2796) );
 wddl_and U2529 ( .A(n2719), .A_n(n2719_n), .B(n2725), .B_n(n2725_n), .Y_n(n3412_n), .Y(n3412) );
 wddl_and U2530 ( .A(n2724), .A_n(n2724_n), .B(n2721), .B_n(n2721_n), .Y_n(n3411_n), .Y(n3411) );
 wddl_and U2531 ( .A(n2675), .A_n(n2675_n), .B(n2552), .B_n(n2552_n), .Y_n(n3306_n), .Y(n3306) );
 wddl_and U2532 ( .A(n2614), .A_n(n2614_n), .B(n2708), .B_n(n2708_n), .Y_n(n3273_n), .Y(n3273) );
 wddl_inv U2533 ( .A(n2724), .A_n(n2724_n), .Y_n(n3380_n), .Y(n3380) );
 wddl_inv U2534 ( .A(n2718), .A_n(n2718_n), .Y_n(n3251_n), .Y(n3251) );
 wddl_inv U2535 ( .A(n2726), .A_n(n2726_n), .Y_n(n3424_n), .Y(n3424) );
endmodule

